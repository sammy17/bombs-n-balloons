`timescale 1ns / 1ps

module block_ram(clk, addr, dout);
	parameter BLOCK_SIZE = 12; // 4 bit R, 4 bit G, 4 bit B
	parameter ADDR_SIZE = 16;
	input clk;
	input [ADDR_SIZE-1:0] addr;
	output reg [BLOCK_SIZE-1:0] dout;

	always @* begin
		case(addr)
			0: dout = 12'h000;
			1: dout = 12'h000;
			2: dout = 12'h000;
			3: dout = 12'h000;
			4: dout = 12'h000;
			5: dout = 12'h000;
			6: dout = 12'h000;
			7: dout = 12'h000;
			8: dout = 12'h000;
			9: dout = 12'h000;
			10: dout = 12'h000;
			11: dout = 12'h000;
			12: dout = 12'h000;
			13: dout = 12'h000;
			14: dout = 12'h000;
			15: dout = 12'h000;
			16: dout = 12'h000;
			17: dout = 12'h000;
			18: dout = 12'h000;
			19: dout = 12'h000;
			20: dout = 12'h000;
			21: dout = 12'h210;
			22: dout = 12'h320;
			23: dout = 12'h320;
			24: dout = 12'h320;
			25: dout = 12'h320;
			26: dout = 12'h320;
			27: dout = 12'h320;
			28: dout = 12'h000;
			29: dout = 12'h000;
			30: dout = 12'h000;
			31: dout = 12'h000;
			32: dout = 12'h000;
			33: dout = 12'h000;
			34: dout = 12'h000;
			35: dout = 12'h000;
			36: dout = 12'h000;
			37: dout = 12'h000;
			38: dout = 12'h000;
			39: dout = 12'h000;

			40: dout = 12'h000;
			41: dout = 12'h000;
			42: dout = 12'h000;
			43: dout = 12'h000;
			44: dout = 12'h000;
			45: dout = 12'h000;
			46: dout = 12'h000;
			47: dout = 12'h000;
			48: dout = 12'h000;
			49: dout = 12'h000;
			50: dout = 12'h000;
			51: dout = 12'h000;
			52: dout = 12'h000;
			53: dout = 12'h000;
			54: dout = 12'h000;
			55: dout = 12'h000;
			56: dout = 12'h000;
			57: dout = 12'h000;
			58: dout = 12'h000;
			59: dout = 12'h000;
			60: dout = 12'h543;
			61: dout = 12'h631;
			62: dout = 12'h631;
			63: dout = 12'h631;
			64: dout = 12'h631;
			65: dout = 12'h631;
			66: dout = 12'h631;
			67: dout = 12'h963;
			68: dout = 12'h321;
			69: dout = 12'h000;
			70: dout = 12'h000;
			71: dout = 12'h000;
			72: dout = 12'h000;
			73: dout = 12'h000;
			74: dout = 12'h000;
			75: dout = 12'h000;
			76: dout = 12'h000;
			77: dout = 12'h000;
			78: dout = 12'h000;
			79: dout = 12'h000;

			80: dout = 12'h000;
			81: dout = 12'h000;
			82: dout = 12'h000;
			83: dout = 12'h000;
			84: dout = 12'h000;
			85: dout = 12'h000;
			86: dout = 12'h000;
			87: dout = 12'h000;
			88: dout = 12'h000;
			89: dout = 12'h000;
			90: dout = 12'h000;
			91: dout = 12'h000;
			92: dout = 12'h000;
			93: dout = 12'h000;
			94: dout = 12'h000;
			95: dout = 12'h000;
			96: dout = 12'h000;
			97: dout = 12'h000;
			98: dout = 12'h000;
			99: dout = 12'h000;
			100: dout = 12'hfc8;
			101: dout = 12'h963;
			102: dout = 12'h752;
			103: dout = 12'h752;
			104: dout = 12'h752;
			105: dout = 12'h752;
			106: dout = 12'h752;
			107: dout = 12'hfc8;
			108: dout = 12'h853;
			109: dout = 12'h210;
			110: dout = 12'h000;
			111: dout = 12'h000;
			112: dout = 12'h000;
			113: dout = 12'h000;
			114: dout = 12'h000;
			115: dout = 12'h000;
			116: dout = 12'h000;
			117: dout = 12'h000;
			118: dout = 12'h000;
			119: dout = 12'h000;

			120: dout = 12'h000;
			121: dout = 12'h000;
			122: dout = 12'h000;
			123: dout = 12'h000;
			124: dout = 12'h000;
			125: dout = 12'h000;
			126: dout = 12'h000;
			127: dout = 12'h000;
			128: dout = 12'h000;
			129: dout = 12'h000;
			130: dout = 12'h000;
			131: dout = 12'h000;
			132: dout = 12'h000;
			133: dout = 12'h000;
			134: dout = 12'h000;
			135: dout = 12'h000;
			136: dout = 12'h000;
			137: dout = 12'h000;
			138: dout = 12'h000;
			139: dout = 12'h000;
			140: dout = 12'hfc8;
			141: dout = 12'hfc8;
			142: dout = 12'hfc8;
			143: dout = 12'hfc8;
			144: dout = 12'hfc8;
			145: dout = 12'hfc8;
			146: dout = 12'hfc8;
			147: dout = 12'hfc8;
			148: dout = 12'h853;
			149: dout = 12'h210;
			150: dout = 12'h000;
			151: dout = 12'h000;
			152: dout = 12'h000;
			153: dout = 12'h000;
			154: dout = 12'h000;
			155: dout = 12'h000;
			156: dout = 12'h000;
			157: dout = 12'h000;
			158: dout = 12'h000;
			159: dout = 12'h000;

			160: dout = 12'h000;
			161: dout = 12'h000;
			162: dout = 12'h000;
			163: dout = 12'h000;
			164: dout = 12'h000;
			165: dout = 12'h000;
			166: dout = 12'h000;
			167: dout = 12'h000;
			168: dout = 12'h000;
			169: dout = 12'h000;
			170: dout = 12'h000;
			171: dout = 12'h000;
			172: dout = 12'h000;
			173: dout = 12'h000;
			174: dout = 12'h000;
			175: dout = 12'h000;
			176: dout = 12'h000;
			177: dout = 12'h000;
			178: dout = 12'h000;
			179: dout = 12'h000;
			180: dout = 12'hfc8;
			181: dout = 12'hfc8;
			182: dout = 12'hfc8;
			183: dout = 12'hfc8;
			184: dout = 12'hfc8;
			185: dout = 12'hfc8;
			186: dout = 12'hfc8;
			187: dout = 12'hfc8;
			188: dout = 12'h853;
			189: dout = 12'h210;
			190: dout = 12'h000;
			191: dout = 12'h000;
			192: dout = 12'h000;
			193: dout = 12'h000;
			194: dout = 12'h000;
			195: dout = 12'h000;
			196: dout = 12'h000;
			197: dout = 12'h000;
			198: dout = 12'h000;
			199: dout = 12'h000;

			200: dout = 12'h000;
			201: dout = 12'h000;
			202: dout = 12'h000;
			203: dout = 12'h000;
			204: dout = 12'h000;
			205: dout = 12'h000;
			206: dout = 12'h000;
			207: dout = 12'h000;
			208: dout = 12'h000;
			209: dout = 12'h000;
			210: dout = 12'h000;
			211: dout = 12'h000;
			212: dout = 12'h000;
			213: dout = 12'h000;
			214: dout = 12'h000;
			215: dout = 12'h000;
			216: dout = 12'h000;
			217: dout = 12'h000;
			218: dout = 12'h000;
			219: dout = 12'h420;
			220: dout = 12'h853;
			221: dout = 12'h432;
			222: dout = 12'hb96;
			223: dout = 12'ha85;
			224: dout = 12'h532;
			225: dout = 12'h853;
			226: dout = 12'h853;
			227: dout = 12'hfc8;
			228: dout = 12'h853;
			229: dout = 12'h210;
			230: dout = 12'h000;
			231: dout = 12'h000;
			232: dout = 12'h000;
			233: dout = 12'h000;
			234: dout = 12'h000;
			235: dout = 12'h000;
			236: dout = 12'h000;
			237: dout = 12'h000;
			238: dout = 12'h000;
			239: dout = 12'h000;

			240: dout = 12'h000;
			241: dout = 12'h000;
			242: dout = 12'h000;
			243: dout = 12'h000;
			244: dout = 12'h000;
			245: dout = 12'h000;
			246: dout = 12'h000;
			247: dout = 12'h000;
			248: dout = 12'h000;
			249: dout = 12'h000;
			250: dout = 12'h000;
			251: dout = 12'h000;
			252: dout = 12'h000;
			253: dout = 12'h000;
			254: dout = 12'h000;
			255: dout = 12'h000;
			256: dout = 12'h000;
			257: dout = 12'h000;
			258: dout = 12'h000;
			259: dout = 12'h210;
			260: dout = 12'h210;
			261: dout = 12'h000;
			262: dout = 12'h432;
			263: dout = 12'h322;
			264: dout = 12'h000;
			265: dout = 12'h210;
			266: dout = 12'h210;
			267: dout = 12'h653;
			268: dout = 12'h321;
			269: dout = 12'h100;
			270: dout = 12'h000;
			271: dout = 12'h000;
			272: dout = 12'h000;
			273: dout = 12'h000;
			274: dout = 12'h000;
			275: dout = 12'h000;
			276: dout = 12'h000;
			277: dout = 12'h000;
			278: dout = 12'h000;
			279: dout = 12'h000;

			280: dout = 12'h000;
			281: dout = 12'h000;
			282: dout = 12'h000;
			283: dout = 12'h000;
			284: dout = 12'h000;
			285: dout = 12'h000;
			286: dout = 12'h000;
			287: dout = 12'h000;
			288: dout = 12'h000;
			289: dout = 12'h000;
			290: dout = 12'h000;
			291: dout = 12'h000;
			292: dout = 12'h000;
			293: dout = 12'h000;
			294: dout = 12'h000;
			295: dout = 12'h000;
			296: dout = 12'h000;
			297: dout = 12'h000;
			298: dout = 12'h100;
			299: dout = 12'h611;
			300: dout = 12'h600;
			301: dout = 12'h622;
			302: dout = 12'h200;
			303: dout = 12'h200;
			304: dout = 12'h611;
			305: dout = 12'h600;
			306: dout = 12'h622;
			307: dout = 12'h000;
			308: dout = 12'h000;
			309: dout = 12'h000;
			310: dout = 12'h000;
			311: dout = 12'h000;
			312: dout = 12'h000;
			313: dout = 12'h000;
			314: dout = 12'h000;
			315: dout = 12'h000;
			316: dout = 12'h000;
			317: dout = 12'h000;
			318: dout = 12'h000;
			319: dout = 12'h000;

			320: dout = 12'h000;
			321: dout = 12'h000;
			322: dout = 12'h000;
			323: dout = 12'h000;
			324: dout = 12'h000;
			325: dout = 12'h000;
			326: dout = 12'h000;
			327: dout = 12'h000;
			328: dout = 12'h000;
			329: dout = 12'h000;
			330: dout = 12'h000;
			331: dout = 12'h000;
			332: dout = 12'h000;
			333: dout = 12'h000;
			334: dout = 12'h000;
			335: dout = 12'h000;
			336: dout = 12'h000;
			337: dout = 12'h000;
			338: dout = 12'h200;
			339: dout = 12'hf35;
			340: dout = 12'hf22;
			341: dout = 12'hf44;
			342: dout = 12'h511;
			343: dout = 12'h712;
			344: dout = 12'hf34;
			345: dout = 12'hf22;
			346: dout = 12'hf55;
			347: dout = 12'h000;
			348: dout = 12'h000;
			349: dout = 12'h000;
			350: dout = 12'h000;
			351: dout = 12'h000;
			352: dout = 12'h000;
			353: dout = 12'h000;
			354: dout = 12'h000;
			355: dout = 12'h000;
			356: dout = 12'h000;
			357: dout = 12'h000;
			358: dout = 12'h000;
			359: dout = 12'h000;

			360: dout = 12'h000;
			361: dout = 12'h000;
			362: dout = 12'h000;
			363: dout = 12'h000;
			364: dout = 12'h000;
			365: dout = 12'h000;
			366: dout = 12'h000;
			367: dout = 12'h000;
			368: dout = 12'h000;
			369: dout = 12'h000;
			370: dout = 12'h000;
			371: dout = 12'h000;
			372: dout = 12'h000;
			373: dout = 12'h000;
			374: dout = 12'h000;
			375: dout = 12'h000;
			376: dout = 12'h000;
			377: dout = 12'h000;
			378: dout = 12'h200;
			379: dout = 12'hf34;
			380: dout = 12'hf34;
			381: dout = 12'hf22;
			382: dout = 12'h500;
			383: dout = 12'h712;
			384: dout = 12'hf34;
			385: dout = 12'hf34;
			386: dout = 12'hf11;
			387: dout = 12'h000;
			388: dout = 12'h000;
			389: dout = 12'h000;
			390: dout = 12'h000;
			391: dout = 12'h000;
			392: dout = 12'h000;
			393: dout = 12'h000;
			394: dout = 12'h000;
			395: dout = 12'h000;
			396: dout = 12'h000;
			397: dout = 12'h000;
			398: dout = 12'h000;
			399: dout = 12'h000;

			400: dout = 12'h000;
			401: dout = 12'h000;
			402: dout = 12'h000;
			403: dout = 12'h000;
			404: dout = 12'h000;
			405: dout = 12'h000;
			406: dout = 12'h000;
			407: dout = 12'h000;
			408: dout = 12'h000;
			409: dout = 12'h000;
			410: dout = 12'h000;
			411: dout = 12'h000;
			412: dout = 12'h000;
			413: dout = 12'h000;
			414: dout = 12'h000;
			415: dout = 12'h000;
			416: dout = 12'h000;
			417: dout = 12'h000;
			418: dout = 12'h000;
			419: dout = 12'h000;
			420: dout = 12'h000;
			421: dout = 12'h000;
			422: dout = 12'h000;
			423: dout = 12'h000;
			424: dout = 12'h000;
			425: dout = 12'h000;
			426: dout = 12'h000;
			427: dout = 12'h000;
			428: dout = 12'h000;
			429: dout = 12'h000;
			430: dout = 12'h000;
			431: dout = 12'h000;
			432: dout = 12'h000;
			433: dout = 12'h000;
			434: dout = 12'h000;
			435: dout = 12'h000;
			436: dout = 12'h000;
			437: dout = 12'h000;
			438: dout = 12'h000;
			439: dout = 12'h000;

			440: dout = 12'h000;
			441: dout = 12'h000;
			442: dout = 12'h333;
			443: dout = 12'h222;
			444: dout = 12'h000;
			445: dout = 12'h000;
			446: dout = 12'h000;
			447: dout = 12'h000;
			448: dout = 12'h000;
			449: dout = 12'h000;
			450: dout = 12'h000;
			451: dout = 12'h000;
			452: dout = 12'h000;
			453: dout = 12'h000;
			454: dout = 12'h000;
			455: dout = 12'h000;
			456: dout = 12'h000;
			457: dout = 12'h000;
			458: dout = 12'h000;
			459: dout = 12'h000;
			460: dout = 12'hda7;
			461: dout = 12'hda7;
			462: dout = 12'hda7;
			463: dout = 12'hda7;
			464: dout = 12'hda7;
			465: dout = 12'hda7;
			466: dout = 12'hda7;
			467: dout = 12'hda7;
			468: dout = 12'h321;
			469: dout = 12'h000;
			470: dout = 12'h000;
			471: dout = 12'h000;
			472: dout = 12'h000;
			473: dout = 12'h000;
			474: dout = 12'h000;
			475: dout = 12'h000;
			476: dout = 12'h000;
			477: dout = 12'h000;
			478: dout = 12'h000;
			479: dout = 12'h000;

			480: dout = 12'h000;
			481: dout = 12'h000;
			482: dout = 12'h555;
			483: dout = 12'h777;
			484: dout = 12'h666;
			485: dout = 12'h666;
			486: dout = 12'h666;
			487: dout = 12'h666;
			488: dout = 12'h666;
			489: dout = 12'h666;
			490: dout = 12'h666;
			491: dout = 12'h444;
			492: dout = 12'h000;
			493: dout = 12'h444;
			494: dout = 12'h000;
			495: dout = 12'h000;
			496: dout = 12'h000;
			497: dout = 12'h000;
			498: dout = 12'h000;
			499: dout = 12'h000;
			500: dout = 12'hfc8;
			501: dout = 12'ha84;
			502: dout = 12'h974;
			503: dout = 12'h974;
			504: dout = 12'hb85;
			505: dout = 12'hfc8;
			506: dout = 12'hfc8;
			507: dout = 12'hfc8;
			508: dout = 12'h332;
			509: dout = 12'h111;
			510: dout = 12'h111;
			511: dout = 12'h000;
			512: dout = 12'h000;
			513: dout = 12'h000;
			514: dout = 12'h000;
			515: dout = 12'h000;
			516: dout = 12'h000;
			517: dout = 12'h000;
			518: dout = 12'h000;
			519: dout = 12'h000;

			520: dout = 12'h000;
			521: dout = 12'h000;
			522: dout = 12'h555;
			523: dout = 12'h888;
			524: dout = 12'h888;
			525: dout = 12'h888;
			526: dout = 12'h888;
			527: dout = 12'h888;
			528: dout = 12'h888;
			529: dout = 12'h999;
			530: dout = 12'h999;
			531: dout = 12'h888;
			532: dout = 12'h444;
			533: dout = 12'h333;
			534: dout = 12'h000;
			535: dout = 12'h000;
			536: dout = 12'h000;
			537: dout = 12'h000;
			538: dout = 12'h000;
			539: dout = 12'h000;
			540: dout = 12'hb85;
			541: dout = 12'ha97;
			542: dout = 12'ha97;
			543: dout = 12'ha97;
			544: dout = 12'ha97;
			545: dout = 12'hc95;
			546: dout = 12'hfc8;
			547: dout = 12'h975;
			548: dout = 12'h211;
			549: dout = 12'h333;
			550: dout = 12'h333;
			551: dout = 12'h000;
			552: dout = 12'h300;
			553: dout = 12'h000;
			554: dout = 12'h000;
			555: dout = 12'h000;
			556: dout = 12'h000;
			557: dout = 12'h000;
			558: dout = 12'h000;
			559: dout = 12'h000;

			560: dout = 12'h000;
			561: dout = 12'h000;
			562: dout = 12'h333;
			563: dout = 12'h555;
			564: dout = 12'h555;
			565: dout = 12'h555;
			566: dout = 12'h555;
			567: dout = 12'h666;
			568: dout = 12'h666;
			569: dout = 12'h777;
			570: dout = 12'h999;
			571: dout = 12'h999;
			572: dout = 12'h999;
			573: dout = 12'h000;
			574: dout = 12'h000;
			575: dout = 12'h100;
			576: dout = 12'h100;
			577: dout = 12'h100;
			578: dout = 12'h100;
			579: dout = 12'h000;
			580: dout = 12'h631;
			581: dout = 12'hedb;
			582: dout = 12'hedc;
			583: dout = 12'hedd;
			584: dout = 12'hdba;
			585: dout = 12'h741;
			586: dout = 12'hb96;
			587: dout = 12'h432;
			588: dout = 12'h000;
			589: dout = 12'h333;
			590: dout = 12'h333;
			591: dout = 12'h100;
			592: dout = 12'h700;
			593: dout = 12'h100;
			594: dout = 12'h000;
			595: dout = 12'h000;
			596: dout = 12'h000;
			597: dout = 12'h000;
			598: dout = 12'h000;
			599: dout = 12'h000;

			600: dout = 12'h000;
			601: dout = 12'h000;
			602: dout = 12'h000;
			603: dout = 12'h000;
			604: dout = 12'h000;
			605: dout = 12'h000;
			606: dout = 12'h000;
			607: dout = 12'h555;
			608: dout = 12'h666;
			609: dout = 12'h666;
			610: dout = 12'h777;
			611: dout = 12'h888;
			612: dout = 12'h888;
			613: dout = 12'h000;
			614: dout = 12'h000;
			615: dout = 12'h500;
			616: dout = 12'h700;
			617: dout = 12'h700;
			618: dout = 12'h600;
			619: dout = 12'h000;
			620: dout = 12'h631;
			621: dout = 12'hda7;
			622: dout = 12'h963;
			623: dout = 12'ha74;
			624: dout = 12'hc96;
			625: dout = 12'h531;
			626: dout = 12'h100;
			627: dout = 12'heb7;
			628: dout = 12'h332;
			629: dout = 12'h333;
			630: dout = 12'h333;
			631: dout = 12'h100;
			632: dout = 12'h700;
			633: dout = 12'h700;
			634: dout = 12'h100;
			635: dout = 12'h000;
			636: dout = 12'h000;
			637: dout = 12'h000;
			638: dout = 12'h000;
			639: dout = 12'h000;

			640: dout = 12'h000;
			641: dout = 12'h000;
			642: dout = 12'h000;
			643: dout = 12'h000;
			644: dout = 12'h000;
			645: dout = 12'h000;
			646: dout = 12'h000;
			647: dout = 12'h000;
			648: dout = 12'h000;
			649: dout = 12'h000;
			650: dout = 12'h000;
			651: dout = 12'h000;
			652: dout = 12'h000;
			653: dout = 12'h000;
			654: dout = 12'h000;
			655: dout = 12'h500;
			656: dout = 12'h300;
			657: dout = 12'h200;
			658: dout = 12'h600;
			659: dout = 12'h000;
			660: dout = 12'h631;
			661: dout = 12'h631;
			662: dout = 12'h631;
			663: dout = 12'h631;
			664: dout = 12'h631;
			665: dout = 12'h742;
			666: dout = 12'hfc8;
			667: dout = 12'h000;
			668: dout = 12'h444;
			669: dout = 12'h555;
			670: dout = 12'h333;
			671: dout = 12'h100;
			672: dout = 12'h700;
			673: dout = 12'h700;
			674: dout = 12'h700;
			675: dout = 12'h200;
			676: dout = 12'h000;
			677: dout = 12'h000;
			678: dout = 12'h000;
			679: dout = 12'h000;

			680: dout = 12'h000;
			681: dout = 12'h000;
			682: dout = 12'h000;
			683: dout = 12'h000;
			684: dout = 12'h000;
			685: dout = 12'h000;
			686: dout = 12'h000;
			687: dout = 12'h000;
			688: dout = 12'h000;
			689: dout = 12'h000;
			690: dout = 12'h111;
			691: dout = 12'h633;
			692: dout = 12'hc00;
			693: dout = 12'hc00;
			694: dout = 12'h100;
			695: dout = 12'h500;
			696: dout = 12'h700;
			697: dout = 12'h400;
			698: dout = 12'h100;
			699: dout = 12'h600;
			700: dout = 12'h000;
			701: dout = 12'h531;
			702: dout = 12'h631;
			703: dout = 12'h631;
			704: dout = 12'h631;
			705: dout = 12'h531;
			706: dout = 12'h211;
			707: dout = 12'h444;
			708: dout = 12'h555;
			709: dout = 12'h222;
			710: dout = 12'h300;
			711: dout = 12'h600;
			712: dout = 12'h700;
			713: dout = 12'h700;
			714: dout = 12'h100;
			715: dout = 12'h000;
			716: dout = 12'h000;
			717: dout = 12'h000;
			718: dout = 12'h000;
			719: dout = 12'h000;

			720: dout = 12'h000;
			721: dout = 12'h000;
			722: dout = 12'h000;
			723: dout = 12'h000;
			724: dout = 12'h000;
			725: dout = 12'h000;
			726: dout = 12'h000;
			727: dout = 12'h000;
			728: dout = 12'h000;
			729: dout = 12'h000;
			730: dout = 12'h222;
			731: dout = 12'h744;
			732: dout = 12'he00;
			733: dout = 12'he00;
			734: dout = 12'h100;
			735: dout = 12'h500;
			736: dout = 12'h700;
			737: dout = 12'h400;
			738: dout = 12'h000;
			739: dout = 12'h200;
			740: dout = 12'h500;
			741: dout = 12'h210;
			742: dout = 12'h210;
			743: dout = 12'h210;
			744: dout = 12'h210;
			745: dout = 12'h210;
			746: dout = 12'h333;
			747: dout = 12'h555;
			748: dout = 12'h222;
			749: dout = 12'h000;
			750: dout = 12'h000;
			751: dout = 12'h200;
			752: dout = 12'h200;
			753: dout = 12'h200;
			754: dout = 12'h400;
			755: dout = 12'h100;
			756: dout = 12'h000;
			757: dout = 12'h000;
			758: dout = 12'h000;
			759: dout = 12'h000;

			760: dout = 12'h000;
			761: dout = 12'h000;
			762: dout = 12'h000;
			763: dout = 12'h000;
			764: dout = 12'h000;
			765: dout = 12'h000;
			766: dout = 12'h000;
			767: dout = 12'h000;
			768: dout = 12'h000;
			769: dout = 12'h000;
			770: dout = 12'h222;
			771: dout = 12'h644;
			772: dout = 12'h922;
			773: dout = 12'h922;
			774: dout = 12'h100;
			775: dout = 12'h200;
			776: dout = 12'h300;
			777: dout = 12'h200;
			778: dout = 12'h000;
			779: dout = 12'h300;
			780: dout = 12'h700;
			781: dout = 12'h700;
			782: dout = 12'h740;
			783: dout = 12'h740;
			784: dout = 12'h720;
			785: dout = 12'h861;
			786: dout = 12'h922;
			787: dout = 12'h922;
			788: dout = 12'h500;
			789: dout = 12'h100;
			790: dout = 12'h100;
			791: dout = 12'h300;
			792: dout = 12'h300;
			793: dout = 12'h300;
			794: dout = 12'h700;
			795: dout = 12'h200;
			796: dout = 12'h000;
			797: dout = 12'h000;
			798: dout = 12'h000;
			799: dout = 12'h000;

			800: dout = 12'h000;
			801: dout = 12'h000;
			802: dout = 12'h000;
			803: dout = 12'h000;
			804: dout = 12'h000;
			805: dout = 12'h000;
			806: dout = 12'h000;
			807: dout = 12'h000;
			808: dout = 12'h000;
			809: dout = 12'h000;
			810: dout = 12'h111;
			811: dout = 12'h333;
			812: dout = 12'h333;
			813: dout = 12'h333;
			814: dout = 12'h000;
			815: dout = 12'h000;
			816: dout = 12'h000;
			817: dout = 12'h000;
			818: dout = 12'h100;
			819: dout = 12'h700;
			820: dout = 12'h700;
			821: dout = 12'hd00;
			822: dout = 12'hf61;
			823: dout = 12'hf71;
			824: dout = 12'hf61;
			825: dout = 12'hf91;
			826: dout = 12'he00;
			827: dout = 12'he00;
			828: dout = 12'h700;
			829: dout = 12'h200;
			830: dout = 12'h200;
			831: dout = 12'h500;
			832: dout = 12'h500;
			833: dout = 12'h500;
			834: dout = 12'h700;
			835: dout = 12'h200;
			836: dout = 12'h000;
			837: dout = 12'h000;
			838: dout = 12'h000;
			839: dout = 12'h000;

			840: dout = 12'h000;
			841: dout = 12'h000;
			842: dout = 12'h000;
			843: dout = 12'h000;
			844: dout = 12'h000;
			845: dout = 12'h000;
			846: dout = 12'h000;
			847: dout = 12'h000;
			848: dout = 12'h000;
			849: dout = 12'h000;
			850: dout = 12'h000;
			851: dout = 12'h000;
			852: dout = 12'h000;
			853: dout = 12'h000;
			854: dout = 12'h000;
			855: dout = 12'h000;
			856: dout = 12'h000;
			857: dout = 12'h000;
			858: dout = 12'h100;
			859: dout = 12'h700;
			860: dout = 12'h700;
			861: dout = 12'hd00;
			862: dout = 12'he10;
			863: dout = 12'hf71;
			864: dout = 12'hfa1;
			865: dout = 12'he10;
			866: dout = 12'he00;
			867: dout = 12'he00;
			868: dout = 12'h300;
			869: dout = 12'h000;
			870: dout = 12'h100;
			871: dout = 12'h100;
			872: dout = 12'h100;
			873: dout = 12'h000;
			874: dout = 12'h600;
			875: dout = 12'h200;
			876: dout = 12'h000;
			877: dout = 12'h000;
			878: dout = 12'h000;
			879: dout = 12'h000;

			880: dout = 12'h000;
			881: dout = 12'h000;
			882: dout = 12'h000;
			883: dout = 12'h000;
			884: dout = 12'h000;
			885: dout = 12'h000;
			886: dout = 12'h000;
			887: dout = 12'h000;
			888: dout = 12'h000;
			889: dout = 12'h000;
			890: dout = 12'h000;
			891: dout = 12'h000;
			892: dout = 12'h000;
			893: dout = 12'h000;
			894: dout = 12'h000;
			895: dout = 12'h000;
			896: dout = 12'h000;
			897: dout = 12'h000;
			898: dout = 12'h100;
			899: dout = 12'h700;
			900: dout = 12'h700;
			901: dout = 12'hd00;
			902: dout = 12'hf91;
			903: dout = 12'hf81;
			904: dout = 12'he40;
			905: dout = 12'hfd1;
			906: dout = 12'he00;
			907: dout = 12'he00;
			908: dout = 12'h300;
			909: dout = 12'h333;
			910: dout = 12'h933;
			911: dout = 12'he00;
			912: dout = 12'hd00;
			913: dout = 12'h000;
			914: dout = 12'h600;
			915: dout = 12'h200;
			916: dout = 12'h000;
			917: dout = 12'h000;
			918: dout = 12'h000;
			919: dout = 12'h000;

			920: dout = 12'h000;
			921: dout = 12'h000;
			922: dout = 12'h000;
			923: dout = 12'h000;
			924: dout = 12'h000;
			925: dout = 12'h000;
			926: dout = 12'h000;
			927: dout = 12'h000;
			928: dout = 12'h000;
			929: dout = 12'h000;
			930: dout = 12'h000;
			931: dout = 12'h000;
			932: dout = 12'h000;
			933: dout = 12'h000;
			934: dout = 12'h000;
			935: dout = 12'h000;
			936: dout = 12'h000;
			937: dout = 12'h000;
			938: dout = 12'h200;
			939: dout = 12'he00;
			940: dout = 12'he00;
			941: dout = 12'h300;
			942: dout = 12'h500;
			943: dout = 12'h800;
			944: dout = 12'h800;
			945: dout = 12'h810;
			946: dout = 12'h800;
			947: dout = 12'h100;
			948: dout = 12'h000;
			949: dout = 12'h333;
			950: dout = 12'h933;
			951: dout = 12'he00;
			952: dout = 12'hd00;
			953: dout = 12'h000;
			954: dout = 12'h000;
			955: dout = 12'h000;
			956: dout = 12'h000;
			957: dout = 12'h000;
			958: dout = 12'h000;
			959: dout = 12'h000;

			960: dout = 12'h000;
			961: dout = 12'h000;
			962: dout = 12'h000;
			963: dout = 12'h000;
			964: dout = 12'h000;
			965: dout = 12'h000;
			966: dout = 12'h000;
			967: dout = 12'h000;
			968: dout = 12'h000;
			969: dout = 12'h000;
			970: dout = 12'h000;
			971: dout = 12'h000;
			972: dout = 12'h000;
			973: dout = 12'h000;
			974: dout = 12'h000;
			975: dout = 12'h000;
			976: dout = 12'h000;
			977: dout = 12'h000;
			978: dout = 12'h200;
			979: dout = 12'he00;
			980: dout = 12'h900;
			981: dout = 12'h600;
			982: dout = 12'h300;
			983: dout = 12'h100;
			984: dout = 12'h100;
			985: dout = 12'h100;
			986: dout = 12'h100;
			987: dout = 12'h500;
			988: dout = 12'h100;
			989: dout = 12'h333;
			990: dout = 12'h644;
			991: dout = 12'h744;
			992: dout = 12'h733;
			993: dout = 12'h000;
			994: dout = 12'h000;
			995: dout = 12'h000;
			996: dout = 12'h000;
			997: dout = 12'h000;
			998: dout = 12'h000;
			999: dout = 12'h000;

			1000: dout = 12'h000;
			1001: dout = 12'h000;
			1002: dout = 12'h000;
			1003: dout = 12'h000;
			1004: dout = 12'h000;
			1005: dout = 12'h000;
			1006: dout = 12'h000;
			1007: dout = 12'h000;
			1008: dout = 12'h000;
			1009: dout = 12'h000;
			1010: dout = 12'h000;
			1011: dout = 12'h000;
			1012: dout = 12'h000;
			1013: dout = 12'h000;
			1014: dout = 12'h000;
			1015: dout = 12'h000;
			1016: dout = 12'h000;
			1017: dout = 12'h000;
			1018: dout = 12'h100;
			1019: dout = 12'ha00;
			1020: dout = 12'h700;
			1021: dout = 12'h700;
			1022: dout = 12'h500;
			1023: dout = 12'h400;
			1024: dout = 12'h400;
			1025: dout = 12'h400;
			1026: dout = 12'h400;
			1027: dout = 12'h700;
			1028: dout = 12'h400;
			1029: dout = 12'h311;
			1030: dout = 12'h222;
			1031: dout = 12'h222;
			1032: dout = 12'h222;
			1033: dout = 12'h000;
			1034: dout = 12'h000;
			1035: dout = 12'h000;
			1036: dout = 12'h000;
			1037: dout = 12'h000;
			1038: dout = 12'h000;
			1039: dout = 12'h000;

			1040: dout = 12'h000;
			1041: dout = 12'h000;
			1042: dout = 12'h000;
			1043: dout = 12'h000;
			1044: dout = 12'h000;
			1045: dout = 12'h000;
			1046: dout = 12'h000;
			1047: dout = 12'h000;
			1048: dout = 12'h000;
			1049: dout = 12'h000;
			1050: dout = 12'h000;
			1051: dout = 12'h000;
			1052: dout = 12'h000;
			1053: dout = 12'h000;
			1054: dout = 12'h000;
			1055: dout = 12'h000;
			1056: dout = 12'h000;
			1057: dout = 12'h000;
			1058: dout = 12'h000;
			1059: dout = 12'h400;
			1060: dout = 12'ha00;
			1061: dout = 12'h500;
			1062: dout = 12'h400;
			1063: dout = 12'h400;
			1064: dout = 12'h400;
			1065: dout = 12'h400;
			1066: dout = 12'h400;
			1067: dout = 12'h400;
			1068: dout = 12'h800;
			1069: dout = 12'h700;
			1070: dout = 12'h300;
			1071: dout = 12'h000;
			1072: dout = 12'h000;
			1073: dout = 12'h000;
			1074: dout = 12'h000;
			1075: dout = 12'h000;
			1076: dout = 12'h000;
			1077: dout = 12'h000;
			1078: dout = 12'h000;
			1079: dout = 12'h000;

			1080: dout = 12'h000;
			1081: dout = 12'h000;
			1082: dout = 12'h000;
			1083: dout = 12'h000;
			1084: dout = 12'h000;
			1085: dout = 12'h000;
			1086: dout = 12'h000;
			1087: dout = 12'h000;
			1088: dout = 12'h000;
			1089: dout = 12'h000;
			1090: dout = 12'h000;
			1091: dout = 12'h000;
			1092: dout = 12'h000;
			1093: dout = 12'h000;
			1094: dout = 12'h000;
			1095: dout = 12'h000;
			1096: dout = 12'h000;
			1097: dout = 12'h000;
			1098: dout = 12'h000;
			1099: dout = 12'h000;
			1100: dout = 12'hc11;
			1101: dout = 12'h400;
			1102: dout = 12'h100;
			1103: dout = 12'h100;
			1104: dout = 12'h100;
			1105: dout = 12'h100;
			1106: dout = 12'h100;
			1107: dout = 12'h000;
			1108: dout = 12'h900;
			1109: dout = 12'hc00;
			1110: dout = 12'h700;
			1111: dout = 12'h000;
			1112: dout = 12'h000;
			1113: dout = 12'h000;
			1114: dout = 12'h000;
			1115: dout = 12'h000;
			1116: dout = 12'h000;
			1117: dout = 12'h000;
			1118: dout = 12'h000;
			1119: dout = 12'h000;

			1120: dout = 12'h000;
			1121: dout = 12'h000;
			1122: dout = 12'h000;
			1123: dout = 12'h000;
			1124: dout = 12'h000;
			1125: dout = 12'h000;
			1126: dout = 12'h000;
			1127: dout = 12'h000;
			1128: dout = 12'h000;
			1129: dout = 12'h000;
			1130: dout = 12'h000;
			1131: dout = 12'h000;
			1132: dout = 12'h000;
			1133: dout = 12'h000;
			1134: dout = 12'h000;
			1135: dout = 12'h000;
			1136: dout = 12'h000;
			1137: dout = 12'h000;
			1138: dout = 12'h000;
			1139: dout = 12'h000;
			1140: dout = 12'h555;
			1141: dout = 12'hc11;
			1142: dout = 12'ha00;
			1143: dout = 12'h700;
			1144: dout = 12'h700;
			1145: dout = 12'h700;
			1146: dout = 12'h700;
			1147: dout = 12'h000;
			1148: dout = 12'h000;
			1149: dout = 12'h000;
			1150: dout = 12'h000;
			1151: dout = 12'h000;
			1152: dout = 12'h000;
			1153: dout = 12'h000;
			1154: dout = 12'h000;
			1155: dout = 12'h000;
			1156: dout = 12'h000;
			1157: dout = 12'h000;
			1158: dout = 12'h000;
			1159: dout = 12'h000;

			1160: dout = 12'h000;
			1161: dout = 12'h000;
			1162: dout = 12'h000;
			1163: dout = 12'h000;
			1164: dout = 12'h000;
			1165: dout = 12'h000;
			1166: dout = 12'h000;
			1167: dout = 12'h000;
			1168: dout = 12'h000;
			1169: dout = 12'h000;
			1170: dout = 12'h000;
			1171: dout = 12'h000;
			1172: dout = 12'h000;
			1173: dout = 12'h000;
			1174: dout = 12'h000;
			1175: dout = 12'h000;
			1176: dout = 12'h000;
			1177: dout = 12'h000;
			1178: dout = 12'h000;
			1179: dout = 12'h000;
			1180: dout = 12'h555;
			1181: dout = 12'hc11;
			1182: dout = 12'ha00;
			1183: dout = 12'h400;
			1184: dout = 12'h200;
			1185: dout = 12'h600;
			1186: dout = 12'h000;
			1187: dout = 12'h600;
			1188: dout = 12'h700;
			1189: dout = 12'hb00;
			1190: dout = 12'h800;
			1191: dout = 12'h000;
			1192: dout = 12'h000;
			1193: dout = 12'h000;
			1194: dout = 12'h000;
			1195: dout = 12'h000;
			1196: dout = 12'h000;
			1197: dout = 12'h000;
			1198: dout = 12'h000;
			1199: dout = 12'h000;

			1200: dout = 12'h000;
			1201: dout = 12'h000;
			1202: dout = 12'h000;
			1203: dout = 12'h000;
			1204: dout = 12'h000;
			1205: dout = 12'h000;
			1206: dout = 12'h000;
			1207: dout = 12'h000;
			1208: dout = 12'h000;
			1209: dout = 12'h000;
			1210: dout = 12'h000;
			1211: dout = 12'h000;
			1212: dout = 12'h000;
			1213: dout = 12'h000;
			1214: dout = 12'h000;
			1215: dout = 12'h000;
			1216: dout = 12'h000;
			1217: dout = 12'h000;
			1218: dout = 12'h200;
			1219: dout = 12'hb00;
			1220: dout = 12'hc11;
			1221: dout = 12'h900;
			1222: dout = 12'h400;
			1223: dout = 12'h000;
			1224: dout = 12'h000;
			1225: dout = 12'h100;
			1226: dout = 12'h000;
			1227: dout = 12'h100;
			1228: dout = 12'ha00;
			1229: dout = 12'hd00;
			1230: dout = 12'h800;
			1231: dout = 12'h000;
			1232: dout = 12'h000;
			1233: dout = 12'h000;
			1234: dout = 12'h000;
			1235: dout = 12'h000;
			1236: dout = 12'h000;
			1237: dout = 12'h000;
			1238: dout = 12'h000;
			1239: dout = 12'h000;

			1240: dout = 12'h000;
			1241: dout = 12'h000;
			1242: dout = 12'h000;
			1243: dout = 12'h000;
			1244: dout = 12'h000;
			1245: dout = 12'h000;
			1246: dout = 12'h000;
			1247: dout = 12'h000;
			1248: dout = 12'h000;
			1249: dout = 12'h000;
			1250: dout = 12'h000;
			1251: dout = 12'h000;
			1252: dout = 12'h000;
			1253: dout = 12'h000;
			1254: dout = 12'h000;
			1255: dout = 12'h000;
			1256: dout = 12'h000;
			1257: dout = 12'h000;
			1258: dout = 12'h100;
			1259: dout = 12'h833;
			1260: dout = 12'he00;
			1261: dout = 12'h800;
			1262: dout = 12'h500;
			1263: dout = 12'h200;
			1264: dout = 12'h000;
			1265: dout = 12'h000;
			1266: dout = 12'h000;
			1267: dout = 12'h400;
			1268: dout = 12'h800;
			1269: dout = 12'h922;
			1270: dout = 12'h522;
			1271: dout = 12'h000;
			1272: dout = 12'h000;
			1273: dout = 12'h000;
			1274: dout = 12'h000;
			1275: dout = 12'h000;
			1276: dout = 12'h000;
			1277: dout = 12'h000;
			1278: dout = 12'h000;
			1279: dout = 12'h000;

			1280: dout = 12'h000;
			1281: dout = 12'h000;
			1282: dout = 12'h000;
			1283: dout = 12'h000;
			1284: dout = 12'h000;
			1285: dout = 12'h000;
			1286: dout = 12'h000;
			1287: dout = 12'h000;
			1288: dout = 12'h000;
			1289: dout = 12'h000;
			1290: dout = 12'h000;
			1291: dout = 12'h000;
			1292: dout = 12'h000;
			1293: dout = 12'h000;
			1294: dout = 12'h000;
			1295: dout = 12'h000;
			1296: dout = 12'h000;
			1297: dout = 12'h000;
			1298: dout = 12'h322;
			1299: dout = 12'h933;
			1300: dout = 12'he00;
			1301: dout = 12'h800;
			1302: dout = 12'h500;
			1303: dout = 12'h200;
			1304: dout = 12'h000;
			1305: dout = 12'h000;
			1306: dout = 12'h000;
			1307: dout = 12'h700;
			1308: dout = 12'h900;
			1309: dout = 12'h922;
			1310: dout = 12'h622;
			1311: dout = 12'h111;
			1312: dout = 12'h000;
			1313: dout = 12'h000;
			1314: dout = 12'h000;
			1315: dout = 12'h000;
			1316: dout = 12'h000;
			1317: dout = 12'h000;
			1318: dout = 12'h000;
			1319: dout = 12'h000;

			1320: dout = 12'h000;
			1321: dout = 12'h000;
			1322: dout = 12'h000;
			1323: dout = 12'h000;
			1324: dout = 12'h000;
			1325: dout = 12'h000;
			1326: dout = 12'h000;
			1327: dout = 12'h000;
			1328: dout = 12'h000;
			1329: dout = 12'h000;
			1330: dout = 12'h000;
			1331: dout = 12'h000;
			1332: dout = 12'h000;
			1333: dout = 12'h000;
			1334: dout = 12'h000;
			1335: dout = 12'h000;
			1336: dout = 12'h000;
			1337: dout = 12'h322;
			1338: dout = 12'h833;
			1339: dout = 12'he00;
			1340: dout = 12'he00;
			1341: dout = 12'ha00;
			1342: dout = 12'h300;
			1343: dout = 12'h000;
			1344: dout = 12'h000;
			1345: dout = 12'h000;
			1346: dout = 12'h000;
			1347: dout = 12'h500;
			1348: dout = 12'hc00;
			1349: dout = 12'he00;
			1350: dout = 12'hb22;
			1351: dout = 12'h633;
			1352: dout = 12'h300;
			1353: dout = 12'h000;
			1354: dout = 12'h000;
			1355: dout = 12'h000;
			1356: dout = 12'h000;
			1357: dout = 12'h000;
			1358: dout = 12'h000;
			1359: dout = 12'h000;

			1360: dout = 12'h000;
			1361: dout = 12'h000;
			1362: dout = 12'h000;
			1363: dout = 12'h000;
			1364: dout = 12'h000;
			1365: dout = 12'h000;
			1366: dout = 12'h000;
			1367: dout = 12'h000;
			1368: dout = 12'h000;
			1369: dout = 12'h000;
			1370: dout = 12'h000;
			1371: dout = 12'h000;
			1372: dout = 12'h000;
			1373: dout = 12'h000;
			1374: dout = 12'h000;
			1375: dout = 12'h000;
			1376: dout = 12'h222;
			1377: dout = 12'h833;
			1378: dout = 12'he00;
			1379: dout = 12'he00;
			1380: dout = 12'he00;
			1381: dout = 12'he00;
			1382: dout = 12'h400;
			1383: dout = 12'h000;
			1384: dout = 12'h000;
			1385: dout = 12'h000;
			1386: dout = 12'h000;
			1387: dout = 12'h000;
			1388: dout = 12'ha00;
			1389: dout = 12'he00;
			1390: dout = 12'he00;
			1391: dout = 12'he00;
			1392: dout = 12'hd00;
			1393: dout = 12'h000;
			1394: dout = 12'h000;
			1395: dout = 12'h000;
			1396: dout = 12'h000;
			1397: dout = 12'h000;
			1398: dout = 12'h000;
			1399: dout = 12'h000;

			1400: dout = 12'h000;
			1401: dout = 12'h000;
			1402: dout = 12'h000;
			1403: dout = 12'h000;
			1404: dout = 12'h000;
			1405: dout = 12'h000;
			1406: dout = 12'h000;
			1407: dout = 12'h000;
			1408: dout = 12'h000;
			1409: dout = 12'h000;
			1410: dout = 12'h000;
			1411: dout = 12'h000;
			1412: dout = 12'h000;
			1413: dout = 12'h000;
			1414: dout = 12'h000;
			1415: dout = 12'h000;
			1416: dout = 12'h222;
			1417: dout = 12'h555;
			1418: dout = 12'h555;
			1419: dout = 12'h555;
			1420: dout = 12'h555;
			1421: dout = 12'h000;
			1422: dout = 12'h000;
			1423: dout = 12'h000;
			1424: dout = 12'h000;
			1425: dout = 12'h000;
			1426: dout = 12'h000;
			1427: dout = 12'h000;
			1428: dout = 12'h444;
			1429: dout = 12'h555;
			1430: dout = 12'h555;
			1431: dout = 12'h555;
			1432: dout = 12'h444;
			1433: dout = 12'h000;
			1434: dout = 12'h000;
			1435: dout = 12'h000;
			1436: dout = 12'h000;
			1437: dout = 12'h000;
			1438: dout = 12'h000;
			1439: dout = 12'h000;

			1440: dout = 12'h000;
			1441: dout = 12'h000;
			1442: dout = 12'h000;
			1443: dout = 12'h000;
			1444: dout = 12'h000;
			1445: dout = 12'h000;
			1446: dout = 12'h000;
			1447: dout = 12'h000;
			1448: dout = 12'h000;
			1449: dout = 12'h000;
			1450: dout = 12'h000;
			1451: dout = 12'h000;
			1452: dout = 12'h000;
			1453: dout = 12'h000;
			1454: dout = 12'h000;
			1455: dout = 12'h000;
			1456: dout = 12'h750;
			1457: dout = 12'hed0;
			1458: dout = 12'hed0;
			1459: dout = 12'hed0;
			1460: dout = 12'hec1;
			1461: dout = 12'h220;
			1462: dout = 12'h000;
			1463: dout = 12'h000;
			1464: dout = 12'h000;
			1465: dout = 12'h000;
			1466: dout = 12'h000;
			1467: dout = 12'h000;
			1468: dout = 12'hc91;
			1469: dout = 12'hed0;
			1470: dout = 12'hed0;
			1471: dout = 12'hed0;
			1472: dout = 12'hd72;
			1473: dout = 12'h000;
			1474: dout = 12'h000;
			1475: dout = 12'h000;
			1476: dout = 12'h000;
			1477: dout = 12'h000;
			1478: dout = 12'h000;
			1479: dout = 12'h000;

			1480: dout = 12'h000;
			1481: dout = 12'h000;
			1482: dout = 12'h000;
			1483: dout = 12'h000;
			1484: dout = 12'h000;
			1485: dout = 12'h000;
			1486: dout = 12'h000;
			1487: dout = 12'h000;
			1488: dout = 12'h000;
			1489: dout = 12'h000;
			1490: dout = 12'h000;
			1491: dout = 12'h000;
			1492: dout = 12'h000;
			1493: dout = 12'h000;
			1494: dout = 12'h000;
			1495: dout = 12'h000;
			1496: dout = 12'h630;
			1497: dout = 12'hfc0;
			1498: dout = 12'hff0;
			1499: dout = 12'hfe0;
			1500: dout = 12'hfa1;
			1501: dout = 12'h210;
			1502: dout = 12'h000;
			1503: dout = 12'h000;
			1504: dout = 12'h000;
			1505: dout = 12'h000;
			1506: dout = 12'h000;
			1507: dout = 12'h000;
			1508: dout = 12'he81;
			1509: dout = 12'hfe0;
			1510: dout = 12'hfe0;
			1511: dout = 12'hfd0;
			1512: dout = 12'hf82;
			1513: dout = 12'h000;
			1514: dout = 12'h000;
			1515: dout = 12'h000;
			1516: dout = 12'h000;
			1517: dout = 12'h000;
			1518: dout = 12'h000;
			1519: dout = 12'h000;

			1520: dout = 12'h000;
			1521: dout = 12'h000;
			1522: dout = 12'h000;
			1523: dout = 12'h000;
			1524: dout = 12'h000;
			1525: dout = 12'h000;
			1526: dout = 12'h000;
			1527: dout = 12'h000;
			1528: dout = 12'h000;
			1529: dout = 12'h000;
			1530: dout = 12'h000;
			1531: dout = 12'h000;
			1532: dout = 12'h000;
			1533: dout = 12'h000;
			1534: dout = 12'h000;
			1535: dout = 12'h000;
			1536: dout = 12'h210;
			1537: dout = 12'hf82;
			1538: dout = 12'hfd0;
			1539: dout = 12'hfc0;
			1540: dout = 12'ha41;
			1541: dout = 12'h210;
			1542: dout = 12'h000;
			1543: dout = 12'h000;
			1544: dout = 12'h000;
			1545: dout = 12'h000;
			1546: dout = 12'h000;
			1547: dout = 12'h000;
			1548: dout = 12'h631;
			1549: dout = 12'hd62;
			1550: dout = 12'hfe0;
			1551: dout = 12'hfd0;
			1552: dout = 12'hd71;
			1553: dout = 12'h000;
			1554: dout = 12'h000;
			1555: dout = 12'h000;
			1556: dout = 12'h000;
			1557: dout = 12'h000;
			1558: dout = 12'h000;
			1559: dout = 12'h000;

			1560: dout = 12'h000;
			1561: dout = 12'h000;
			1562: dout = 12'h000;
			1563: dout = 12'h000;
			1564: dout = 12'h000;
			1565: dout = 12'h000;
			1566: dout = 12'h000;
			1567: dout = 12'h000;
			1568: dout = 12'h000;
			1569: dout = 12'h000;
			1570: dout = 12'h000;
			1571: dout = 12'h000;
			1572: dout = 12'h000;
			1573: dout = 12'h000;
			1574: dout = 12'h000;
			1575: dout = 12'h000;
			1576: dout = 12'h000;
			1577: dout = 12'h841;
			1578: dout = 12'hf92;
			1579: dout = 12'hfc0;
			1580: dout = 12'h000;
			1581: dout = 12'h000;
			1582: dout = 12'h000;
			1583: dout = 12'h000;
			1584: dout = 12'h000;
			1585: dout = 12'h000;
			1586: dout = 12'h000;
			1587: dout = 12'h000;
			1588: dout = 12'h000;
			1589: dout = 12'h941;
			1590: dout = 12'hfc1;
			1591: dout = 12'hcb0;
			1592: dout = 12'h420;
			1593: dout = 12'h000;
			1594: dout = 12'h000;
			1595: dout = 12'h000;
			1596: dout = 12'h000;
			1597: dout = 12'h000;
			1598: dout = 12'h000;
			1599: dout = 12'h000;

			1600: dout = 12'h000;
			1601: dout = 12'h000;
			1602: dout = 12'h000;
			1603: dout = 12'h000;
			1604: dout = 12'h000;
			1605: dout = 12'h000;
			1606: dout = 12'h000;
			1607: dout = 12'h000;
			1608: dout = 12'h000;
			1609: dout = 12'h000;
			1610: dout = 12'h000;
			1611: dout = 12'h000;
			1612: dout = 12'h000;
			1613: dout = 12'h000;
			1614: dout = 12'h000;
			1615: dout = 12'h000;
			1616: dout = 12'h000;
			1617: dout = 12'h000;
			1618: dout = 12'ha51;
			1619: dout = 12'hea1;
			1620: dout = 12'h000;
			1621: dout = 12'h000;
			1622: dout = 12'h000;
			1623: dout = 12'h000;
			1624: dout = 12'h000;
			1625: dout = 12'h000;
			1626: dout = 12'h000;
			1627: dout = 12'h000;
			1628: dout = 12'h210;
			1629: dout = 12'h941;
			1630: dout = 12'h530;
			1631: dout = 12'h220;
			1632: dout = 12'h000;
			1633: dout = 12'h000;
			1634: dout = 12'h000;
			1635: dout = 12'h000;
			1636: dout = 12'h000;
			1637: dout = 12'h000;
			1638: dout = 12'h000;
			1639: dout = 12'h000;

			1640: dout = 12'h000;
			1641: dout = 12'h000;
			1642: dout = 12'h000;
			1643: dout = 12'h000;
			1644: dout = 12'h000;
			1645: dout = 12'h000;
			1646: dout = 12'h000;
			1647: dout = 12'h000;
			1648: dout = 12'h000;
			1649: dout = 12'h000;
			1650: dout = 12'h000;
			1651: dout = 12'h000;
			1652: dout = 12'h000;
			1653: dout = 12'h000;
			1654: dout = 12'h000;
			1655: dout = 12'h000;
			1656: dout = 12'h000;
			1657: dout = 12'h000;
			1658: dout = 12'h000;
			1659: dout = 12'h520;
			1660: dout = 12'h000;
			1661: dout = 12'h000;
			1662: dout = 12'h000;
			1663: dout = 12'h000;
			1664: dout = 12'h000;
			1665: dout = 12'h000;
			1666: dout = 12'h000;
			1667: dout = 12'h000;
			1668: dout = 12'h000;
			1669: dout = 12'h210;
			1670: dout = 12'h841;
			1671: dout = 12'h000;
			1672: dout = 12'h000;
			1673: dout = 12'h000;
			1674: dout = 12'h000;
			1675: dout = 12'h000;
			1676: dout = 12'h000;
			1677: dout = 12'h000;
			1678: dout = 12'h000;
			1679: dout = 12'h000;

			1680: dout = 12'h000;
			1681: dout = 12'h000;
			1682: dout = 12'h000;
			1683: dout = 12'h000;
			1684: dout = 12'h000;
			1685: dout = 12'h000;
			1686: dout = 12'h000;
			1687: dout = 12'h000;
			1688: dout = 12'h000;
			1689: dout = 12'h000;
			1690: dout = 12'h000;
			1691: dout = 12'h000;
			1692: dout = 12'h000;
			1693: dout = 12'h000;
			1694: dout = 12'h000;
			1695: dout = 12'h000;
			1696: dout = 12'h000;
			1697: dout = 12'h000;
			1698: dout = 12'h000;
			1699: dout = 12'h210;
			1700: dout = 12'h000;
			1701: dout = 12'h000;
			1702: dout = 12'h000;
			1703: dout = 12'h000;
			1704: dout = 12'h000;
			1705: dout = 12'h000;
			1706: dout = 12'h000;
			1707: dout = 12'h000;
			1708: dout = 12'h000;
			1709: dout = 12'h000;
			1710: dout = 12'h000;
			1711: dout = 12'h000;
			1712: dout = 12'h000;
			1713: dout = 12'h000;
			1714: dout = 12'h000;
			1715: dout = 12'h000;
			1716: dout = 12'h000;
			1717: dout = 12'h000;
			1718: dout = 12'h000;
			1719: dout = 12'h000;

			1720: dout = 12'h000;
			1721: dout = 12'h000;
			1722: dout = 12'h000;
			1723: dout = 12'h000;
			1724: dout = 12'h000;
			1725: dout = 12'h000;
			1726: dout = 12'h000;
			1727: dout = 12'h000;
			1728: dout = 12'h000;
			1729: dout = 12'h000;
			1730: dout = 12'h000;
			1731: dout = 12'h000;
			1732: dout = 12'h000;
			1733: dout = 12'h000;
			1734: dout = 12'h000;
			1735: dout = 12'h000;
			1736: dout = 12'h000;
			1737: dout = 12'h000;
			1738: dout = 12'h000;
			1739: dout = 12'h000;
			1740: dout = 12'h000;
			1741: dout = 12'h000;
			1742: dout = 12'h000;
			1743: dout = 12'h000;
			1744: dout = 12'h000;
			1745: dout = 12'h000;
			1746: dout = 12'h000;
			1747: dout = 12'h000;
			1748: dout = 12'h000;
			1749: dout = 12'h000;
			1750: dout = 12'h000;
			1751: dout = 12'h000;
			1752: dout = 12'h000;
			1753: dout = 12'h000;
			1754: dout = 12'h000;
			1755: dout = 12'h000;
			1756: dout = 12'h000;
			1757: dout = 12'h000;
			1758: dout = 12'h000;
			1759: dout = 12'h000;

			1760: dout = 12'h000;
			1761: dout = 12'h000;
			1762: dout = 12'h000;
			1763: dout = 12'h000;
			1764: dout = 12'h000;
			1765: dout = 12'h000;
			1766: dout = 12'h000;
			1767: dout = 12'h000;
			1768: dout = 12'h000;
			1769: dout = 12'h000;
			1770: dout = 12'h000;
			1771: dout = 12'h000;
			1772: dout = 12'h000;
			1773: dout = 12'h000;
			1774: dout = 12'h000;
			1775: dout = 12'h000;
			1776: dout = 12'h000;
			1777: dout = 12'h000;
			1778: dout = 12'h000;
			1779: dout = 12'h000;
			1780: dout = 12'h000;
			1781: dout = 12'h210;
			1782: dout = 12'h320;
			1783: dout = 12'h320;
			1784: dout = 12'h320;
			1785: dout = 12'h320;
			1786: dout = 12'h320;
			1787: dout = 12'h320;
			1788: dout = 12'h000;
			1789: dout = 12'h000;
			1790: dout = 12'h000;
			1791: dout = 12'h000;
			1792: dout = 12'h000;
			1793: dout = 12'h000;
			1794: dout = 12'h000;
			1795: dout = 12'h000;
			1796: dout = 12'h000;
			1797: dout = 12'h000;
			1798: dout = 12'h000;
			1799: dout = 12'h000;

			1800: dout = 12'h000;
			1801: dout = 12'h000;
			1802: dout = 12'h000;
			1803: dout = 12'h000;
			1804: dout = 12'h000;
			1805: dout = 12'h000;
			1806: dout = 12'h000;
			1807: dout = 12'h000;
			1808: dout = 12'h000;
			1809: dout = 12'h000;
			1810: dout = 12'h000;
			1811: dout = 12'h000;
			1812: dout = 12'h000;
			1813: dout = 12'h000;
			1814: dout = 12'h000;
			1815: dout = 12'h000;
			1816: dout = 12'h000;
			1817: dout = 12'h000;
			1818: dout = 12'h000;
			1819: dout = 12'h000;
			1820: dout = 12'h543;
			1821: dout = 12'h631;
			1822: dout = 12'h631;
			1823: dout = 12'h631;
			1824: dout = 12'h631;
			1825: dout = 12'h631;
			1826: dout = 12'h631;
			1827: dout = 12'h963;
			1828: dout = 12'h321;
			1829: dout = 12'h000;
			1830: dout = 12'h000;
			1831: dout = 12'h000;
			1832: dout = 12'h000;
			1833: dout = 12'h000;
			1834: dout = 12'h000;
			1835: dout = 12'h000;
			1836: dout = 12'h000;
			1837: dout = 12'h000;
			1838: dout = 12'h000;
			1839: dout = 12'h000;

			1840: dout = 12'h000;
			1841: dout = 12'h000;
			1842: dout = 12'h000;
			1843: dout = 12'h000;
			1844: dout = 12'h000;
			1845: dout = 12'h000;
			1846: dout = 12'h000;
			1847: dout = 12'h000;
			1848: dout = 12'h000;
			1849: dout = 12'h000;
			1850: dout = 12'h000;
			1851: dout = 12'h000;
			1852: dout = 12'h000;
			1853: dout = 12'h000;
			1854: dout = 12'h000;
			1855: dout = 12'h000;
			1856: dout = 12'h000;
			1857: dout = 12'h000;
			1858: dout = 12'h000;
			1859: dout = 12'h000;
			1860: dout = 12'hfc8;
			1861: dout = 12'h963;
			1862: dout = 12'h752;
			1863: dout = 12'h752;
			1864: dout = 12'h752;
			1865: dout = 12'h752;
			1866: dout = 12'h752;
			1867: dout = 12'hfc8;
			1868: dout = 12'h853;
			1869: dout = 12'h210;
			1870: dout = 12'h000;
			1871: dout = 12'h000;
			1872: dout = 12'h000;
			1873: dout = 12'h000;
			1874: dout = 12'h000;
			1875: dout = 12'h000;
			1876: dout = 12'h000;
			1877: dout = 12'h000;
			1878: dout = 12'h000;
			1879: dout = 12'h000;

			1880: dout = 12'h000;
			1881: dout = 12'h000;
			1882: dout = 12'h000;
			1883: dout = 12'h000;
			1884: dout = 12'h000;
			1885: dout = 12'h000;
			1886: dout = 12'h000;
			1887: dout = 12'h000;
			1888: dout = 12'h000;
			1889: dout = 12'h000;
			1890: dout = 12'h000;
			1891: dout = 12'h000;
			1892: dout = 12'h000;
			1893: dout = 12'h000;
			1894: dout = 12'h000;
			1895: dout = 12'h000;
			1896: dout = 12'h000;
			1897: dout = 12'h000;
			1898: dout = 12'h000;
			1899: dout = 12'h000;
			1900: dout = 12'hfc8;
			1901: dout = 12'hfc8;
			1902: dout = 12'hfc8;
			1903: dout = 12'hfc8;
			1904: dout = 12'hfc8;
			1905: dout = 12'hfc8;
			1906: dout = 12'hfc8;
			1907: dout = 12'hfc8;
			1908: dout = 12'h853;
			1909: dout = 12'h210;
			1910: dout = 12'h000;
			1911: dout = 12'h000;
			1912: dout = 12'h000;
			1913: dout = 12'h000;
			1914: dout = 12'h000;
			1915: dout = 12'h000;
			1916: dout = 12'h000;
			1917: dout = 12'h000;
			1918: dout = 12'h000;
			1919: dout = 12'h000;

			1920: dout = 12'h000;
			1921: dout = 12'h000;
			1922: dout = 12'h000;
			1923: dout = 12'h000;
			1924: dout = 12'h000;
			1925: dout = 12'h000;
			1926: dout = 12'h000;
			1927: dout = 12'h000;
			1928: dout = 12'h000;
			1929: dout = 12'h000;
			1930: dout = 12'h000;
			1931: dout = 12'h000;
			1932: dout = 12'h000;
			1933: dout = 12'h000;
			1934: dout = 12'h000;
			1935: dout = 12'h000;
			1936: dout = 12'h000;
			1937: dout = 12'h000;
			1938: dout = 12'h000;
			1939: dout = 12'h000;
			1940: dout = 12'hfc8;
			1941: dout = 12'hfc8;
			1942: dout = 12'hfc8;
			1943: dout = 12'hfc8;
			1944: dout = 12'hfc8;
			1945: dout = 12'hfc8;
			1946: dout = 12'hfc8;
			1947: dout = 12'hfc8;
			1948: dout = 12'h853;
			1949: dout = 12'h210;
			1950: dout = 12'h000;
			1951: dout = 12'h000;
			1952: dout = 12'h000;
			1953: dout = 12'h000;
			1954: dout = 12'h000;
			1955: dout = 12'h000;
			1956: dout = 12'h000;
			1957: dout = 12'h000;
			1958: dout = 12'h000;
			1959: dout = 12'h000;

			1960: dout = 12'h000;
			1961: dout = 12'h000;
			1962: dout = 12'h000;
			1963: dout = 12'h000;
			1964: dout = 12'h000;
			1965: dout = 12'h000;
			1966: dout = 12'h000;
			1967: dout = 12'h000;
			1968: dout = 12'h000;
			1969: dout = 12'h000;
			1970: dout = 12'h000;
			1971: dout = 12'h000;
			1972: dout = 12'h000;
			1973: dout = 12'h000;
			1974: dout = 12'h000;
			1975: dout = 12'h000;
			1976: dout = 12'h000;
			1977: dout = 12'h000;
			1978: dout = 12'h000;
			1979: dout = 12'h420;
			1980: dout = 12'h853;
			1981: dout = 12'h432;
			1982: dout = 12'hb96;
			1983: dout = 12'ha85;
			1984: dout = 12'h532;
			1985: dout = 12'h853;
			1986: dout = 12'h853;
			1987: dout = 12'hfc8;
			1988: dout = 12'h853;
			1989: dout = 12'h210;
			1990: dout = 12'h000;
			1991: dout = 12'h000;
			1992: dout = 12'h000;
			1993: dout = 12'h000;
			1994: dout = 12'h000;
			1995: dout = 12'h000;
			1996: dout = 12'h000;
			1997: dout = 12'h000;
			1998: dout = 12'h000;
			1999: dout = 12'h000;

			2000: dout = 12'h000;
			2001: dout = 12'h000;
			2002: dout = 12'h000;
			2003: dout = 12'h000;
			2004: dout = 12'h000;
			2005: dout = 12'h000;
			2006: dout = 12'h000;
			2007: dout = 12'h000;
			2008: dout = 12'h000;
			2009: dout = 12'h000;
			2010: dout = 12'h000;
			2011: dout = 12'h000;
			2012: dout = 12'h000;
			2013: dout = 12'h000;
			2014: dout = 12'h000;
			2015: dout = 12'h000;
			2016: dout = 12'h000;
			2017: dout = 12'h000;
			2018: dout = 12'h000;
			2019: dout = 12'h210;
			2020: dout = 12'h210;
			2021: dout = 12'h000;
			2022: dout = 12'h432;
			2023: dout = 12'h322;
			2024: dout = 12'h000;
			2025: dout = 12'h210;
			2026: dout = 12'h210;
			2027: dout = 12'h653;
			2028: dout = 12'h321;
			2029: dout = 12'h100;
			2030: dout = 12'h000;
			2031: dout = 12'h000;
			2032: dout = 12'h000;
			2033: dout = 12'h000;
			2034: dout = 12'h000;
			2035: dout = 12'h000;
			2036: dout = 12'h000;
			2037: dout = 12'h000;
			2038: dout = 12'h000;
			2039: dout = 12'h000;

			2040: dout = 12'h000;
			2041: dout = 12'h000;
			2042: dout = 12'h000;
			2043: dout = 12'h000;
			2044: dout = 12'h000;
			2045: dout = 12'h000;
			2046: dout = 12'h000;
			2047: dout = 12'h000;
			2048: dout = 12'h000;
			2049: dout = 12'h000;
			2050: dout = 12'h000;
			2051: dout = 12'h000;
			2052: dout = 12'h000;
			2053: dout = 12'h000;
			2054: dout = 12'h000;
			2055: dout = 12'h000;
			2056: dout = 12'h000;
			2057: dout = 12'h000;
			2058: dout = 12'h100;
			2059: dout = 12'h611;
			2060: dout = 12'h600;
			2061: dout = 12'h622;
			2062: dout = 12'h200;
			2063: dout = 12'h200;
			2064: dout = 12'h611;
			2065: dout = 12'h600;
			2066: dout = 12'h622;
			2067: dout = 12'h000;
			2068: dout = 12'h000;
			2069: dout = 12'h000;
			2070: dout = 12'h000;
			2071: dout = 12'h000;
			2072: dout = 12'h000;
			2073: dout = 12'h000;
			2074: dout = 12'h000;
			2075: dout = 12'h000;
			2076: dout = 12'h000;
			2077: dout = 12'h000;
			2078: dout = 12'h000;
			2079: dout = 12'h000;

			2080: dout = 12'h000;
			2081: dout = 12'h000;
			2082: dout = 12'h000;
			2083: dout = 12'h000;
			2084: dout = 12'h000;
			2085: dout = 12'h000;
			2086: dout = 12'h000;
			2087: dout = 12'h000;
			2088: dout = 12'h000;
			2089: dout = 12'h000;
			2090: dout = 12'h000;
			2091: dout = 12'h000;
			2092: dout = 12'h000;
			2093: dout = 12'h000;
			2094: dout = 12'h000;
			2095: dout = 12'h000;
			2096: dout = 12'h000;
			2097: dout = 12'h000;
			2098: dout = 12'h200;
			2099: dout = 12'hf35;
			2100: dout = 12'hf22;
			2101: dout = 12'hf44;
			2102: dout = 12'h511;
			2103: dout = 12'h712;
			2104: dout = 12'hf34;
			2105: dout = 12'hf22;
			2106: dout = 12'hf55;
			2107: dout = 12'h000;
			2108: dout = 12'h000;
			2109: dout = 12'h000;
			2110: dout = 12'h000;
			2111: dout = 12'h000;
			2112: dout = 12'h000;
			2113: dout = 12'h000;
			2114: dout = 12'h000;
			2115: dout = 12'h000;
			2116: dout = 12'h000;
			2117: dout = 12'h000;
			2118: dout = 12'h000;
			2119: dout = 12'h000;

			2120: dout = 12'h000;
			2121: dout = 12'h000;
			2122: dout = 12'h000;
			2123: dout = 12'h000;
			2124: dout = 12'h000;
			2125: dout = 12'h000;
			2126: dout = 12'h000;
			2127: dout = 12'h000;
			2128: dout = 12'h000;
			2129: dout = 12'h000;
			2130: dout = 12'h000;
			2131: dout = 12'h000;
			2132: dout = 12'h000;
			2133: dout = 12'h000;
			2134: dout = 12'h000;
			2135: dout = 12'h000;
			2136: dout = 12'h000;
			2137: dout = 12'h000;
			2138: dout = 12'h200;
			2139: dout = 12'hf34;
			2140: dout = 12'hf34;
			2141: dout = 12'hf22;
			2142: dout = 12'h500;
			2143: dout = 12'h712;
			2144: dout = 12'hf34;
			2145: dout = 12'hf34;
			2146: dout = 12'hf11;
			2147: dout = 12'h000;
			2148: dout = 12'h000;
			2149: dout = 12'h000;
			2150: dout = 12'h000;
			2151: dout = 12'h000;
			2152: dout = 12'h000;
			2153: dout = 12'h000;
			2154: dout = 12'h000;
			2155: dout = 12'h000;
			2156: dout = 12'h000;
			2157: dout = 12'h000;
			2158: dout = 12'h000;
			2159: dout = 12'h000;

			2160: dout = 12'h000;
			2161: dout = 12'h000;
			2162: dout = 12'h000;
			2163: dout = 12'h000;
			2164: dout = 12'h000;
			2165: dout = 12'h000;
			2166: dout = 12'h000;
			2167: dout = 12'h000;
			2168: dout = 12'h000;
			2169: dout = 12'h000;
			2170: dout = 12'h000;
			2171: dout = 12'h000;
			2172: dout = 12'h000;
			2173: dout = 12'h000;
			2174: dout = 12'h000;
			2175: dout = 12'h000;
			2176: dout = 12'h000;
			2177: dout = 12'h000;
			2178: dout = 12'h000;
			2179: dout = 12'h000;
			2180: dout = 12'h000;
			2181: dout = 12'h000;
			2182: dout = 12'h000;
			2183: dout = 12'h000;
			2184: dout = 12'h000;
			2185: dout = 12'h000;
			2186: dout = 12'h000;
			2187: dout = 12'h000;
			2188: dout = 12'h000;
			2189: dout = 12'h000;
			2190: dout = 12'h000;
			2191: dout = 12'h000;
			2192: dout = 12'h000;
			2193: dout = 12'h000;
			2194: dout = 12'h000;
			2195: dout = 12'h000;
			2196: dout = 12'h000;
			2197: dout = 12'h000;
			2198: dout = 12'h000;
			2199: dout = 12'h000;

			2200: dout = 12'h000;
			2201: dout = 12'h000;
			2202: dout = 12'h333;
			2203: dout = 12'h222;
			2204: dout = 12'h000;
			2205: dout = 12'h000;
			2206: dout = 12'h000;
			2207: dout = 12'h000;
			2208: dout = 12'h000;
			2209: dout = 12'h000;
			2210: dout = 12'h000;
			2211: dout = 12'h000;
			2212: dout = 12'h000;
			2213: dout = 12'h000;
			2214: dout = 12'h000;
			2215: dout = 12'h000;
			2216: dout = 12'h000;
			2217: dout = 12'h000;
			2218: dout = 12'h000;
			2219: dout = 12'h000;
			2220: dout = 12'hda7;
			2221: dout = 12'hda7;
			2222: dout = 12'hda7;
			2223: dout = 12'hda7;
			2224: dout = 12'hda7;
			2225: dout = 12'hda7;
			2226: dout = 12'hda7;
			2227: dout = 12'hda7;
			2228: dout = 12'h321;
			2229: dout = 12'h000;
			2230: dout = 12'h000;
			2231: dout = 12'h000;
			2232: dout = 12'h000;
			2233: dout = 12'h000;
			2234: dout = 12'h000;
			2235: dout = 12'h000;
			2236: dout = 12'h000;
			2237: dout = 12'h000;
			2238: dout = 12'h000;
			2239: dout = 12'h000;

			2240: dout = 12'h000;
			2241: dout = 12'h000;
			2242: dout = 12'h555;
			2243: dout = 12'h777;
			2244: dout = 12'h666;
			2245: dout = 12'h666;
			2246: dout = 12'h666;
			2247: dout = 12'h666;
			2248: dout = 12'h666;
			2249: dout = 12'h666;
			2250: dout = 12'h666;
			2251: dout = 12'h444;
			2252: dout = 12'h000;
			2253: dout = 12'h444;
			2254: dout = 12'h000;
			2255: dout = 12'h000;
			2256: dout = 12'h000;
			2257: dout = 12'h000;
			2258: dout = 12'h000;
			2259: dout = 12'h000;
			2260: dout = 12'hfc8;
			2261: dout = 12'ha84;
			2262: dout = 12'h974;
			2263: dout = 12'h974;
			2264: dout = 12'hb85;
			2265: dout = 12'hfc8;
			2266: dout = 12'hfc8;
			2267: dout = 12'hfc8;
			2268: dout = 12'h332;
			2269: dout = 12'h111;
			2270: dout = 12'h111;
			2271: dout = 12'h000;
			2272: dout = 12'h000;
			2273: dout = 12'h000;
			2274: dout = 12'h000;
			2275: dout = 12'h000;
			2276: dout = 12'h000;
			2277: dout = 12'h000;
			2278: dout = 12'h000;
			2279: dout = 12'h000;

			2280: dout = 12'h000;
			2281: dout = 12'h000;
			2282: dout = 12'h555;
			2283: dout = 12'h888;
			2284: dout = 12'h888;
			2285: dout = 12'h888;
			2286: dout = 12'h888;
			2287: dout = 12'h888;
			2288: dout = 12'h888;
			2289: dout = 12'h999;
			2290: dout = 12'h999;
			2291: dout = 12'h888;
			2292: dout = 12'h444;
			2293: dout = 12'h333;
			2294: dout = 12'h000;
			2295: dout = 12'h000;
			2296: dout = 12'h000;
			2297: dout = 12'h000;
			2298: dout = 12'h000;
			2299: dout = 12'h000;
			2300: dout = 12'hb85;
			2301: dout = 12'ha97;
			2302: dout = 12'ha97;
			2303: dout = 12'ha97;
			2304: dout = 12'ha97;
			2305: dout = 12'hc95;
			2306: dout = 12'hfc8;
			2307: dout = 12'h975;
			2308: dout = 12'h211;
			2309: dout = 12'h333;
			2310: dout = 12'h333;
			2311: dout = 12'h000;
			2312: dout = 12'h300;
			2313: dout = 12'h000;
			2314: dout = 12'h000;
			2315: dout = 12'h000;
			2316: dout = 12'h000;
			2317: dout = 12'h000;
			2318: dout = 12'h000;
			2319: dout = 12'h000;

			2320: dout = 12'h000;
			2321: dout = 12'h000;
			2322: dout = 12'h333;
			2323: dout = 12'h555;
			2324: dout = 12'h555;
			2325: dout = 12'h555;
			2326: dout = 12'h555;
			2327: dout = 12'h666;
			2328: dout = 12'h666;
			2329: dout = 12'h777;
			2330: dout = 12'h999;
			2331: dout = 12'h999;
			2332: dout = 12'h999;
			2333: dout = 12'h000;
			2334: dout = 12'h000;
			2335: dout = 12'h100;
			2336: dout = 12'h100;
			2337: dout = 12'h100;
			2338: dout = 12'h100;
			2339: dout = 12'h000;
			2340: dout = 12'h631;
			2341: dout = 12'hedb;
			2342: dout = 12'hedc;
			2343: dout = 12'hedd;
			2344: dout = 12'hdba;
			2345: dout = 12'h741;
			2346: dout = 12'hb96;
			2347: dout = 12'h432;
			2348: dout = 12'h000;
			2349: dout = 12'h333;
			2350: dout = 12'h333;
			2351: dout = 12'h100;
			2352: dout = 12'h700;
			2353: dout = 12'h100;
			2354: dout = 12'h000;
			2355: dout = 12'h000;
			2356: dout = 12'h000;
			2357: dout = 12'h000;
			2358: dout = 12'h000;
			2359: dout = 12'h000;

			2360: dout = 12'h000;
			2361: dout = 12'h000;
			2362: dout = 12'h000;
			2363: dout = 12'h000;
			2364: dout = 12'h000;
			2365: dout = 12'h000;
			2366: dout = 12'h000;
			2367: dout = 12'h555;
			2368: dout = 12'h666;
			2369: dout = 12'h666;
			2370: dout = 12'h777;
			2371: dout = 12'h888;
			2372: dout = 12'h888;
			2373: dout = 12'h000;
			2374: dout = 12'h000;
			2375: dout = 12'h500;
			2376: dout = 12'h700;
			2377: dout = 12'h700;
			2378: dout = 12'h600;
			2379: dout = 12'h000;
			2380: dout = 12'h631;
			2381: dout = 12'hda7;
			2382: dout = 12'h963;
			2383: dout = 12'ha74;
			2384: dout = 12'hc96;
			2385: dout = 12'h531;
			2386: dout = 12'h100;
			2387: dout = 12'heb7;
			2388: dout = 12'h332;
			2389: dout = 12'h333;
			2390: dout = 12'h333;
			2391: dout = 12'h100;
			2392: dout = 12'h700;
			2393: dout = 12'h700;
			2394: dout = 12'h100;
			2395: dout = 12'h000;
			2396: dout = 12'h000;
			2397: dout = 12'h000;
			2398: dout = 12'h000;
			2399: dout = 12'h000;

			2400: dout = 12'h000;
			2401: dout = 12'h000;
			2402: dout = 12'h000;
			2403: dout = 12'h000;
			2404: dout = 12'h000;
			2405: dout = 12'h000;
			2406: dout = 12'h000;
			2407: dout = 12'h000;
			2408: dout = 12'h000;
			2409: dout = 12'h000;
			2410: dout = 12'h000;
			2411: dout = 12'h000;
			2412: dout = 12'h000;
			2413: dout = 12'h000;
			2414: dout = 12'h000;
			2415: dout = 12'h500;
			2416: dout = 12'h300;
			2417: dout = 12'h200;
			2418: dout = 12'h600;
			2419: dout = 12'h000;
			2420: dout = 12'h631;
			2421: dout = 12'h631;
			2422: dout = 12'h631;
			2423: dout = 12'h631;
			2424: dout = 12'h631;
			2425: dout = 12'h742;
			2426: dout = 12'hfc8;
			2427: dout = 12'h000;
			2428: dout = 12'h444;
			2429: dout = 12'h555;
			2430: dout = 12'h333;
			2431: dout = 12'h100;
			2432: dout = 12'h700;
			2433: dout = 12'h700;
			2434: dout = 12'h700;
			2435: dout = 12'h200;
			2436: dout = 12'h000;
			2437: dout = 12'h000;
			2438: dout = 12'h000;
			2439: dout = 12'h000;

			2440: dout = 12'h000;
			2441: dout = 12'h000;
			2442: dout = 12'h000;
			2443: dout = 12'h000;
			2444: dout = 12'h000;
			2445: dout = 12'h000;
			2446: dout = 12'h000;
			2447: dout = 12'h000;
			2448: dout = 12'h000;
			2449: dout = 12'h000;
			2450: dout = 12'h111;
			2451: dout = 12'h633;
			2452: dout = 12'hc00;
			2453: dout = 12'hc00;
			2454: dout = 12'h100;
			2455: dout = 12'h500;
			2456: dout = 12'h700;
			2457: dout = 12'h400;
			2458: dout = 12'h100;
			2459: dout = 12'h600;
			2460: dout = 12'h000;
			2461: dout = 12'h531;
			2462: dout = 12'h631;
			2463: dout = 12'h631;
			2464: dout = 12'h631;
			2465: dout = 12'h531;
			2466: dout = 12'h211;
			2467: dout = 12'h444;
			2468: dout = 12'h555;
			2469: dout = 12'h222;
			2470: dout = 12'h300;
			2471: dout = 12'h600;
			2472: dout = 12'h700;
			2473: dout = 12'h700;
			2474: dout = 12'h100;
			2475: dout = 12'h000;
			2476: dout = 12'h000;
			2477: dout = 12'h000;
			2478: dout = 12'h000;
			2479: dout = 12'h000;

			2480: dout = 12'h000;
			2481: dout = 12'h000;
			2482: dout = 12'h000;
			2483: dout = 12'h000;
			2484: dout = 12'h000;
			2485: dout = 12'h000;
			2486: dout = 12'h000;
			2487: dout = 12'h000;
			2488: dout = 12'h000;
			2489: dout = 12'h000;
			2490: dout = 12'h222;
			2491: dout = 12'h744;
			2492: dout = 12'he00;
			2493: dout = 12'he00;
			2494: dout = 12'h100;
			2495: dout = 12'h500;
			2496: dout = 12'h700;
			2497: dout = 12'h400;
			2498: dout = 12'h000;
			2499: dout = 12'h200;
			2500: dout = 12'h500;
			2501: dout = 12'h210;
			2502: dout = 12'h210;
			2503: dout = 12'h210;
			2504: dout = 12'h210;
			2505: dout = 12'h210;
			2506: dout = 12'h333;
			2507: dout = 12'h555;
			2508: dout = 12'h222;
			2509: dout = 12'h000;
			2510: dout = 12'h000;
			2511: dout = 12'h200;
			2512: dout = 12'h200;
			2513: dout = 12'h200;
			2514: dout = 12'h400;
			2515: dout = 12'h100;
			2516: dout = 12'h000;
			2517: dout = 12'h000;
			2518: dout = 12'h000;
			2519: dout = 12'h000;

			2520: dout = 12'h000;
			2521: dout = 12'h000;
			2522: dout = 12'h000;
			2523: dout = 12'h000;
			2524: dout = 12'h000;
			2525: dout = 12'h000;
			2526: dout = 12'h000;
			2527: dout = 12'h000;
			2528: dout = 12'h000;
			2529: dout = 12'h000;
			2530: dout = 12'h222;
			2531: dout = 12'h644;
			2532: dout = 12'h922;
			2533: dout = 12'h922;
			2534: dout = 12'h100;
			2535: dout = 12'h200;
			2536: dout = 12'h300;
			2537: dout = 12'h200;
			2538: dout = 12'h000;
			2539: dout = 12'h300;
			2540: dout = 12'h700;
			2541: dout = 12'h700;
			2542: dout = 12'h740;
			2543: dout = 12'h740;
			2544: dout = 12'h720;
			2545: dout = 12'h861;
			2546: dout = 12'h922;
			2547: dout = 12'h922;
			2548: dout = 12'h500;
			2549: dout = 12'h100;
			2550: dout = 12'h100;
			2551: dout = 12'h300;
			2552: dout = 12'h300;
			2553: dout = 12'h300;
			2554: dout = 12'h700;
			2555: dout = 12'h200;
			2556: dout = 12'h000;
			2557: dout = 12'h000;
			2558: dout = 12'h000;
			2559: dout = 12'h000;

			2560: dout = 12'h000;
			2561: dout = 12'h000;
			2562: dout = 12'h000;
			2563: dout = 12'h000;
			2564: dout = 12'h000;
			2565: dout = 12'h000;
			2566: dout = 12'h000;
			2567: dout = 12'h000;
			2568: dout = 12'h000;
			2569: dout = 12'h000;
			2570: dout = 12'h111;
			2571: dout = 12'h333;
			2572: dout = 12'h333;
			2573: dout = 12'h333;
			2574: dout = 12'h000;
			2575: dout = 12'h000;
			2576: dout = 12'h000;
			2577: dout = 12'h000;
			2578: dout = 12'h100;
			2579: dout = 12'h700;
			2580: dout = 12'h700;
			2581: dout = 12'hd00;
			2582: dout = 12'hf61;
			2583: dout = 12'hf71;
			2584: dout = 12'hf61;
			2585: dout = 12'hf91;
			2586: dout = 12'he00;
			2587: dout = 12'he00;
			2588: dout = 12'h700;
			2589: dout = 12'h200;
			2590: dout = 12'h200;
			2591: dout = 12'h500;
			2592: dout = 12'h500;
			2593: dout = 12'h500;
			2594: dout = 12'h700;
			2595: dout = 12'h200;
			2596: dout = 12'h000;
			2597: dout = 12'h000;
			2598: dout = 12'h000;
			2599: dout = 12'h000;

			2600: dout = 12'h000;
			2601: dout = 12'h000;
			2602: dout = 12'h000;
			2603: dout = 12'h000;
			2604: dout = 12'h000;
			2605: dout = 12'h000;
			2606: dout = 12'h000;
			2607: dout = 12'h000;
			2608: dout = 12'h000;
			2609: dout = 12'h000;
			2610: dout = 12'h000;
			2611: dout = 12'h000;
			2612: dout = 12'h000;
			2613: dout = 12'h000;
			2614: dout = 12'h000;
			2615: dout = 12'h000;
			2616: dout = 12'h000;
			2617: dout = 12'h000;
			2618: dout = 12'h100;
			2619: dout = 12'h700;
			2620: dout = 12'h700;
			2621: dout = 12'hd00;
			2622: dout = 12'he10;
			2623: dout = 12'hf71;
			2624: dout = 12'hfa1;
			2625: dout = 12'he10;
			2626: dout = 12'he00;
			2627: dout = 12'he00;
			2628: dout = 12'h300;
			2629: dout = 12'h000;
			2630: dout = 12'h100;
			2631: dout = 12'h100;
			2632: dout = 12'h100;
			2633: dout = 12'h000;
			2634: dout = 12'h600;
			2635: dout = 12'h200;
			2636: dout = 12'h000;
			2637: dout = 12'h000;
			2638: dout = 12'h000;
			2639: dout = 12'h000;

			2640: dout = 12'h000;
			2641: dout = 12'h000;
			2642: dout = 12'h000;
			2643: dout = 12'h000;
			2644: dout = 12'h000;
			2645: dout = 12'h000;
			2646: dout = 12'h000;
			2647: dout = 12'h000;
			2648: dout = 12'h000;
			2649: dout = 12'h000;
			2650: dout = 12'h000;
			2651: dout = 12'h000;
			2652: dout = 12'h000;
			2653: dout = 12'h000;
			2654: dout = 12'h000;
			2655: dout = 12'h000;
			2656: dout = 12'h000;
			2657: dout = 12'h000;
			2658: dout = 12'h100;
			2659: dout = 12'h700;
			2660: dout = 12'h700;
			2661: dout = 12'hd00;
			2662: dout = 12'hf91;
			2663: dout = 12'hf81;
			2664: dout = 12'he40;
			2665: dout = 12'hfd1;
			2666: dout = 12'he00;
			2667: dout = 12'he00;
			2668: dout = 12'h300;
			2669: dout = 12'h333;
			2670: dout = 12'h933;
			2671: dout = 12'he00;
			2672: dout = 12'hd00;
			2673: dout = 12'h000;
			2674: dout = 12'h600;
			2675: dout = 12'h200;
			2676: dout = 12'h000;
			2677: dout = 12'h000;
			2678: dout = 12'h000;
			2679: dout = 12'h000;

			2680: dout = 12'h000;
			2681: dout = 12'h000;
			2682: dout = 12'h000;
			2683: dout = 12'h000;
			2684: dout = 12'h000;
			2685: dout = 12'h000;
			2686: dout = 12'h000;
			2687: dout = 12'h000;
			2688: dout = 12'h000;
			2689: dout = 12'h000;
			2690: dout = 12'h000;
			2691: dout = 12'h000;
			2692: dout = 12'h000;
			2693: dout = 12'h000;
			2694: dout = 12'h000;
			2695: dout = 12'h000;
			2696: dout = 12'h000;
			2697: dout = 12'h000;
			2698: dout = 12'h200;
			2699: dout = 12'he00;
			2700: dout = 12'he00;
			2701: dout = 12'h300;
			2702: dout = 12'h500;
			2703: dout = 12'h800;
			2704: dout = 12'h800;
			2705: dout = 12'h810;
			2706: dout = 12'h800;
			2707: dout = 12'h100;
			2708: dout = 12'h000;
			2709: dout = 12'h333;
			2710: dout = 12'h933;
			2711: dout = 12'he00;
			2712: dout = 12'hd00;
			2713: dout = 12'h000;
			2714: dout = 12'h000;
			2715: dout = 12'h000;
			2716: dout = 12'h000;
			2717: dout = 12'h000;
			2718: dout = 12'h000;
			2719: dout = 12'h000;

			2720: dout = 12'h000;
			2721: dout = 12'h000;
			2722: dout = 12'h000;
			2723: dout = 12'h000;
			2724: dout = 12'h000;
			2725: dout = 12'h000;
			2726: dout = 12'h000;
			2727: dout = 12'h000;
			2728: dout = 12'h000;
			2729: dout = 12'h000;
			2730: dout = 12'h000;
			2731: dout = 12'h000;
			2732: dout = 12'h000;
			2733: dout = 12'h000;
			2734: dout = 12'h000;
			2735: dout = 12'h000;
			2736: dout = 12'h000;
			2737: dout = 12'h000;
			2738: dout = 12'h200;
			2739: dout = 12'he00;
			2740: dout = 12'h900;
			2741: dout = 12'h600;
			2742: dout = 12'h300;
			2743: dout = 12'h100;
			2744: dout = 12'h100;
			2745: dout = 12'h100;
			2746: dout = 12'h100;
			2747: dout = 12'h500;
			2748: dout = 12'h100;
			2749: dout = 12'h333;
			2750: dout = 12'h644;
			2751: dout = 12'h744;
			2752: dout = 12'h733;
			2753: dout = 12'h000;
			2754: dout = 12'h000;
			2755: dout = 12'h000;
			2756: dout = 12'h000;
			2757: dout = 12'h000;
			2758: dout = 12'h000;
			2759: dout = 12'h000;

			2760: dout = 12'h000;
			2761: dout = 12'h000;
			2762: dout = 12'h000;
			2763: dout = 12'h000;
			2764: dout = 12'h000;
			2765: dout = 12'h000;
			2766: dout = 12'h000;
			2767: dout = 12'h000;
			2768: dout = 12'h000;
			2769: dout = 12'h000;
			2770: dout = 12'h000;
			2771: dout = 12'h000;
			2772: dout = 12'h000;
			2773: dout = 12'h000;
			2774: dout = 12'h000;
			2775: dout = 12'h000;
			2776: dout = 12'h000;
			2777: dout = 12'h000;
			2778: dout = 12'h100;
			2779: dout = 12'ha00;
			2780: dout = 12'h700;
			2781: dout = 12'h700;
			2782: dout = 12'h500;
			2783: dout = 12'h400;
			2784: dout = 12'h400;
			2785: dout = 12'h400;
			2786: dout = 12'h400;
			2787: dout = 12'h700;
			2788: dout = 12'h400;
			2789: dout = 12'h311;
			2790: dout = 12'h222;
			2791: dout = 12'h222;
			2792: dout = 12'h222;
			2793: dout = 12'h000;
			2794: dout = 12'h000;
			2795: dout = 12'h000;
			2796: dout = 12'h000;
			2797: dout = 12'h000;
			2798: dout = 12'h000;
			2799: dout = 12'h000;

			2800: dout = 12'h000;
			2801: dout = 12'h000;
			2802: dout = 12'h000;
			2803: dout = 12'h000;
			2804: dout = 12'h000;
			2805: dout = 12'h000;
			2806: dout = 12'h000;
			2807: dout = 12'h000;
			2808: dout = 12'h000;
			2809: dout = 12'h000;
			2810: dout = 12'h000;
			2811: dout = 12'h000;
			2812: dout = 12'h000;
			2813: dout = 12'h000;
			2814: dout = 12'h000;
			2815: dout = 12'h000;
			2816: dout = 12'h000;
			2817: dout = 12'h000;
			2818: dout = 12'h000;
			2819: dout = 12'h400;
			2820: dout = 12'ha00;
			2821: dout = 12'h500;
			2822: dout = 12'h400;
			2823: dout = 12'h400;
			2824: dout = 12'h400;
			2825: dout = 12'h400;
			2826: dout = 12'h400;
			2827: dout = 12'h400;
			2828: dout = 12'h800;
			2829: dout = 12'h700;
			2830: dout = 12'h300;
			2831: dout = 12'h000;
			2832: dout = 12'h000;
			2833: dout = 12'h000;
			2834: dout = 12'h000;
			2835: dout = 12'h000;
			2836: dout = 12'h000;
			2837: dout = 12'h000;
			2838: dout = 12'h000;
			2839: dout = 12'h000;

			2840: dout = 12'h000;
			2841: dout = 12'h000;
			2842: dout = 12'h000;
			2843: dout = 12'h000;
			2844: dout = 12'h000;
			2845: dout = 12'h000;
			2846: dout = 12'h000;
			2847: dout = 12'h000;
			2848: dout = 12'h000;
			2849: dout = 12'h000;
			2850: dout = 12'h000;
			2851: dout = 12'h000;
			2852: dout = 12'h000;
			2853: dout = 12'h000;
			2854: dout = 12'h000;
			2855: dout = 12'h000;
			2856: dout = 12'h000;
			2857: dout = 12'h000;
			2858: dout = 12'h000;
			2859: dout = 12'h000;
			2860: dout = 12'hc11;
			2861: dout = 12'h400;
			2862: dout = 12'h100;
			2863: dout = 12'h100;
			2864: dout = 12'h100;
			2865: dout = 12'h100;
			2866: dout = 12'h100;
			2867: dout = 12'h000;
			2868: dout = 12'h900;
			2869: dout = 12'hc00;
			2870: dout = 12'h700;
			2871: dout = 12'h000;
			2872: dout = 12'h000;
			2873: dout = 12'h000;
			2874: dout = 12'h000;
			2875: dout = 12'h000;
			2876: dout = 12'h000;
			2877: dout = 12'h000;
			2878: dout = 12'h000;
			2879: dout = 12'h000;

			2880: dout = 12'h000;
			2881: dout = 12'h000;
			2882: dout = 12'h000;
			2883: dout = 12'h000;
			2884: dout = 12'h000;
			2885: dout = 12'h000;
			2886: dout = 12'h000;
			2887: dout = 12'h000;
			2888: dout = 12'h000;
			2889: dout = 12'h000;
			2890: dout = 12'h000;
			2891: dout = 12'h000;
			2892: dout = 12'h000;
			2893: dout = 12'h000;
			2894: dout = 12'h000;
			2895: dout = 12'h000;
			2896: dout = 12'h000;
			2897: dout = 12'h000;
			2898: dout = 12'h000;
			2899: dout = 12'h000;
			2900: dout = 12'h555;
			2901: dout = 12'hc11;
			2902: dout = 12'ha00;
			2903: dout = 12'h700;
			2904: dout = 12'h700;
			2905: dout = 12'h700;
			2906: dout = 12'h700;
			2907: dout = 12'h000;
			2908: dout = 12'h000;
			2909: dout = 12'h000;
			2910: dout = 12'h000;
			2911: dout = 12'h000;
			2912: dout = 12'h000;
			2913: dout = 12'h000;
			2914: dout = 12'h000;
			2915: dout = 12'h000;
			2916: dout = 12'h000;
			2917: dout = 12'h000;
			2918: dout = 12'h000;
			2919: dout = 12'h000;

			2920: dout = 12'h000;
			2921: dout = 12'h000;
			2922: dout = 12'h000;
			2923: dout = 12'h000;
			2924: dout = 12'h000;
			2925: dout = 12'h000;
			2926: dout = 12'h000;
			2927: dout = 12'h000;
			2928: dout = 12'h000;
			2929: dout = 12'h000;
			2930: dout = 12'h000;
			2931: dout = 12'h000;
			2932: dout = 12'h000;
			2933: dout = 12'h000;
			2934: dout = 12'h000;
			2935: dout = 12'h000;
			2936: dout = 12'h000;
			2937: dout = 12'h000;
			2938: dout = 12'h000;
			2939: dout = 12'h000;
			2940: dout = 12'h555;
			2941: dout = 12'hc11;
			2942: dout = 12'ha00;
			2943: dout = 12'h400;
			2944: dout = 12'h200;
			2945: dout = 12'h600;
			2946: dout = 12'h000;
			2947: dout = 12'h600;
			2948: dout = 12'h700;
			2949: dout = 12'hb00;
			2950: dout = 12'h800;
			2951: dout = 12'h000;
			2952: dout = 12'h000;
			2953: dout = 12'h000;
			2954: dout = 12'h000;
			2955: dout = 12'h000;
			2956: dout = 12'h000;
			2957: dout = 12'h000;
			2958: dout = 12'h000;
			2959: dout = 12'h000;

			2960: dout = 12'h000;
			2961: dout = 12'h000;
			2962: dout = 12'h000;
			2963: dout = 12'h000;
			2964: dout = 12'h000;
			2965: dout = 12'h000;
			2966: dout = 12'h000;
			2967: dout = 12'h000;
			2968: dout = 12'h000;
			2969: dout = 12'h000;
			2970: dout = 12'h000;
			2971: dout = 12'h000;
			2972: dout = 12'h000;
			2973: dout = 12'h000;
			2974: dout = 12'h000;
			2975: dout = 12'h000;
			2976: dout = 12'h000;
			2977: dout = 12'h000;
			2978: dout = 12'h200;
			2979: dout = 12'hb00;
			2980: dout = 12'hc11;
			2981: dout = 12'h900;
			2982: dout = 12'h400;
			2983: dout = 12'h000;
			2984: dout = 12'h000;
			2985: dout = 12'h100;
			2986: dout = 12'h000;
			2987: dout = 12'h100;
			2988: dout = 12'ha00;
			2989: dout = 12'hd00;
			2990: dout = 12'h800;
			2991: dout = 12'h000;
			2992: dout = 12'h000;
			2993: dout = 12'h000;
			2994: dout = 12'h000;
			2995: dout = 12'h000;
			2996: dout = 12'h000;
			2997: dout = 12'h000;
			2998: dout = 12'h000;
			2999: dout = 12'h000;

			3000: dout = 12'h000;
			3001: dout = 12'h000;
			3002: dout = 12'h000;
			3003: dout = 12'h000;
			3004: dout = 12'h000;
			3005: dout = 12'h000;
			3006: dout = 12'h000;
			3007: dout = 12'h000;
			3008: dout = 12'h000;
			3009: dout = 12'h000;
			3010: dout = 12'h000;
			3011: dout = 12'h000;
			3012: dout = 12'h000;
			3013: dout = 12'h000;
			3014: dout = 12'h000;
			3015: dout = 12'h000;
			3016: dout = 12'h000;
			3017: dout = 12'h000;
			3018: dout = 12'h100;
			3019: dout = 12'h833;
			3020: dout = 12'he00;
			3021: dout = 12'h800;
			3022: dout = 12'h500;
			3023: dout = 12'h200;
			3024: dout = 12'h000;
			3025: dout = 12'h000;
			3026: dout = 12'h000;
			3027: dout = 12'h400;
			3028: dout = 12'h800;
			3029: dout = 12'h922;
			3030: dout = 12'h522;
			3031: dout = 12'h000;
			3032: dout = 12'h000;
			3033: dout = 12'h000;
			3034: dout = 12'h000;
			3035: dout = 12'h000;
			3036: dout = 12'h000;
			3037: dout = 12'h000;
			3038: dout = 12'h000;
			3039: dout = 12'h000;

			3040: dout = 12'h000;
			3041: dout = 12'h000;
			3042: dout = 12'h000;
			3043: dout = 12'h000;
			3044: dout = 12'h000;
			3045: dout = 12'h000;
			3046: dout = 12'h000;
			3047: dout = 12'h000;
			3048: dout = 12'h000;
			3049: dout = 12'h000;
			3050: dout = 12'h000;
			3051: dout = 12'h000;
			3052: dout = 12'h000;
			3053: dout = 12'h000;
			3054: dout = 12'h000;
			3055: dout = 12'h000;
			3056: dout = 12'h000;
			3057: dout = 12'h000;
			3058: dout = 12'h322;
			3059: dout = 12'h933;
			3060: dout = 12'he00;
			3061: dout = 12'h800;
			3062: dout = 12'h500;
			3063: dout = 12'h200;
			3064: dout = 12'h000;
			3065: dout = 12'h000;
			3066: dout = 12'h000;
			3067: dout = 12'h700;
			3068: dout = 12'h900;
			3069: dout = 12'h922;
			3070: dout = 12'h622;
			3071: dout = 12'h111;
			3072: dout = 12'h000;
			3073: dout = 12'h000;
			3074: dout = 12'h000;
			3075: dout = 12'h000;
			3076: dout = 12'h000;
			3077: dout = 12'h000;
			3078: dout = 12'h000;
			3079: dout = 12'h000;

			3080: dout = 12'h000;
			3081: dout = 12'h000;
			3082: dout = 12'h000;
			3083: dout = 12'h000;
			3084: dout = 12'h000;
			3085: dout = 12'h000;
			3086: dout = 12'h000;
			3087: dout = 12'h000;
			3088: dout = 12'h000;
			3089: dout = 12'h000;
			3090: dout = 12'h000;
			3091: dout = 12'h000;
			3092: dout = 12'h000;
			3093: dout = 12'h000;
			3094: dout = 12'h000;
			3095: dout = 12'h000;
			3096: dout = 12'h000;
			3097: dout = 12'h322;
			3098: dout = 12'h833;
			3099: dout = 12'he00;
			3100: dout = 12'he00;
			3101: dout = 12'ha00;
			3102: dout = 12'h300;
			3103: dout = 12'h000;
			3104: dout = 12'h000;
			3105: dout = 12'h000;
			3106: dout = 12'h000;
			3107: dout = 12'h500;
			3108: dout = 12'hc00;
			3109: dout = 12'he00;
			3110: dout = 12'hb22;
			3111: dout = 12'h633;
			3112: dout = 12'h300;
			3113: dout = 12'h000;
			3114: dout = 12'h000;
			3115: dout = 12'h000;
			3116: dout = 12'h000;
			3117: dout = 12'h000;
			3118: dout = 12'h000;
			3119: dout = 12'h000;

			3120: dout = 12'h000;
			3121: dout = 12'h000;
			3122: dout = 12'h000;
			3123: dout = 12'h000;
			3124: dout = 12'h000;
			3125: dout = 12'h000;
			3126: dout = 12'h000;
			3127: dout = 12'h000;
			3128: dout = 12'h000;
			3129: dout = 12'h000;
			3130: dout = 12'h000;
			3131: dout = 12'h000;
			3132: dout = 12'h000;
			3133: dout = 12'h000;
			3134: dout = 12'h000;
			3135: dout = 12'h000;
			3136: dout = 12'h222;
			3137: dout = 12'h833;
			3138: dout = 12'he00;
			3139: dout = 12'he00;
			3140: dout = 12'he00;
			3141: dout = 12'he00;
			3142: dout = 12'h400;
			3143: dout = 12'h000;
			3144: dout = 12'h000;
			3145: dout = 12'h000;
			3146: dout = 12'h000;
			3147: dout = 12'h000;
			3148: dout = 12'ha00;
			3149: dout = 12'he00;
			3150: dout = 12'he00;
			3151: dout = 12'he00;
			3152: dout = 12'hd00;
			3153: dout = 12'h000;
			3154: dout = 12'h000;
			3155: dout = 12'h000;
			3156: dout = 12'h000;
			3157: dout = 12'h000;
			3158: dout = 12'h000;
			3159: dout = 12'h000;

			3160: dout = 12'h000;
			3161: dout = 12'h000;
			3162: dout = 12'h000;
			3163: dout = 12'h000;
			3164: dout = 12'h000;
			3165: dout = 12'h000;
			3166: dout = 12'h000;
			3167: dout = 12'h000;
			3168: dout = 12'h000;
			3169: dout = 12'h000;
			3170: dout = 12'h000;
			3171: dout = 12'h000;
			3172: dout = 12'h000;
			3173: dout = 12'h000;
			3174: dout = 12'h000;
			3175: dout = 12'h000;
			3176: dout = 12'h222;
			3177: dout = 12'h555;
			3178: dout = 12'h555;
			3179: dout = 12'h555;
			3180: dout = 12'h555;
			3181: dout = 12'h000;
			3182: dout = 12'h000;
			3183: dout = 12'h000;
			3184: dout = 12'h000;
			3185: dout = 12'h000;
			3186: dout = 12'h000;
			3187: dout = 12'h000;
			3188: dout = 12'h444;
			3189: dout = 12'h555;
			3190: dout = 12'h555;
			3191: dout = 12'h555;
			3192: dout = 12'h444;
			3193: dout = 12'h000;
			3194: dout = 12'h000;
			3195: dout = 12'h000;
			3196: dout = 12'h000;
			3197: dout = 12'h000;
			3198: dout = 12'h000;
			3199: dout = 12'h000;

			3200: dout = 12'h000;
			3201: dout = 12'h000;
			3202: dout = 12'h000;
			3203: dout = 12'h000;
			3204: dout = 12'h000;
			3205: dout = 12'h000;
			3206: dout = 12'h000;
			3207: dout = 12'h000;
			3208: dout = 12'h000;
			3209: dout = 12'h000;
			3210: dout = 12'h000;
			3211: dout = 12'h000;
			3212: dout = 12'h000;
			3213: dout = 12'h000;
			3214: dout = 12'h000;
			3215: dout = 12'h000;
			3216: dout = 12'h760;
			3217: dout = 12'hed0;
			3218: dout = 12'hed0;
			3219: dout = 12'hed0;
			3220: dout = 12'hec1;
			3221: dout = 12'h420;
			3222: dout = 12'h000;
			3223: dout = 12'h000;
			3224: dout = 12'h000;
			3225: dout = 12'h000;
			3226: dout = 12'h000;
			3227: dout = 12'h000;
			3228: dout = 12'ha81;
			3229: dout = 12'hed0;
			3230: dout = 12'hed0;
			3231: dout = 12'hed0;
			3232: dout = 12'hda1;
			3233: dout = 12'h000;
			3234: dout = 12'h000;
			3235: dout = 12'h000;
			3236: dout = 12'h000;
			3237: dout = 12'h000;
			3238: dout = 12'h000;
			3239: dout = 12'h000;

			3240: dout = 12'h000;
			3241: dout = 12'h000;
			3242: dout = 12'h000;
			3243: dout = 12'h000;
			3244: dout = 12'h000;
			3245: dout = 12'h000;
			3246: dout = 12'h000;
			3247: dout = 12'h000;
			3248: dout = 12'h000;
			3249: dout = 12'h000;
			3250: dout = 12'h000;
			3251: dout = 12'h000;
			3252: dout = 12'h000;
			3253: dout = 12'h000;
			3254: dout = 12'h000;
			3255: dout = 12'h000;
			3256: dout = 12'h750;
			3257: dout = 12'hfd0;
			3258: dout = 12'hfe0;
			3259: dout = 12'hfd0;
			3260: dout = 12'hfa1;
			3261: dout = 12'h941;
			3262: dout = 12'h000;
			3263: dout = 12'h000;
			3264: dout = 12'h000;
			3265: dout = 12'h000;
			3266: dout = 12'h000;
			3267: dout = 12'h000;
			3268: dout = 12'hc81;
			3269: dout = 12'hfe0;
			3270: dout = 12'hfe0;
			3271: dout = 12'hfd0;
			3272: dout = 12'hf82;
			3273: dout = 12'h310;
			3274: dout = 12'h000;
			3275: dout = 12'h000;
			3276: dout = 12'h000;
			3277: dout = 12'h000;
			3278: dout = 12'h000;
			3279: dout = 12'h000;

			3280: dout = 12'h000;
			3281: dout = 12'h000;
			3282: dout = 12'h000;
			3283: dout = 12'h000;
			3284: dout = 12'h000;
			3285: dout = 12'h000;
			3286: dout = 12'h000;
			3287: dout = 12'h000;
			3288: dout = 12'h000;
			3289: dout = 12'h000;
			3290: dout = 12'h000;
			3291: dout = 12'h000;
			3292: dout = 12'h000;
			3293: dout = 12'h000;
			3294: dout = 12'h000;
			3295: dout = 12'h000;
			3296: dout = 12'h000;
			3297: dout = 12'hf91;
			3298: dout = 12'hfe0;
			3299: dout = 12'hfd0;
			3300: dout = 12'hfa1;
			3301: dout = 12'h210;
			3302: dout = 12'h000;
			3303: dout = 12'h000;
			3304: dout = 12'h000;
			3305: dout = 12'h000;
			3306: dout = 12'h000;
			3307: dout = 12'h000;
			3308: dout = 12'h630;
			3309: dout = 12'hfa1;
			3310: dout = 12'hfb1;
			3311: dout = 12'hfa1;
			3312: dout = 12'hf82;
			3313: dout = 12'h210;
			3314: dout = 12'h000;
			3315: dout = 12'h000;
			3316: dout = 12'h000;
			3317: dout = 12'h000;
			3318: dout = 12'h000;
			3319: dout = 12'h000;

			3320: dout = 12'h000;
			3321: dout = 12'h000;
			3322: dout = 12'h000;
			3323: dout = 12'h000;
			3324: dout = 12'h000;
			3325: dout = 12'h000;
			3326: dout = 12'h000;
			3327: dout = 12'h000;
			3328: dout = 12'h000;
			3329: dout = 12'h000;
			3330: dout = 12'h000;
			3331: dout = 12'h000;
			3332: dout = 12'h000;
			3333: dout = 12'h000;
			3334: dout = 12'h000;
			3335: dout = 12'h000;
			3336: dout = 12'h000;
			3337: dout = 12'hfa1;
			3338: dout = 12'hfc0;
			3339: dout = 12'hfa1;
			3340: dout = 12'hfc1;
			3341: dout = 12'h210;
			3342: dout = 12'h000;
			3343: dout = 12'h000;
			3344: dout = 12'h000;
			3345: dout = 12'h000;
			3346: dout = 12'h000;
			3347: dout = 12'h000;
			3348: dout = 12'h000;
			3349: dout = 12'h841;
			3350: dout = 12'hf82;
			3351: dout = 12'hd72;
			3352: dout = 12'hd62;
			3353: dout = 12'h000;
			3354: dout = 12'h000;
			3355: dout = 12'h000;
			3356: dout = 12'h000;
			3357: dout = 12'h000;
			3358: dout = 12'h000;
			3359: dout = 12'h000;

			3360: dout = 12'h000;
			3361: dout = 12'h000;
			3362: dout = 12'h000;
			3363: dout = 12'h000;
			3364: dout = 12'h000;
			3365: dout = 12'h000;
			3366: dout = 12'h000;
			3367: dout = 12'h000;
			3368: dout = 12'h000;
			3369: dout = 12'h000;
			3370: dout = 12'h000;
			3371: dout = 12'h000;
			3372: dout = 12'h000;
			3373: dout = 12'h000;
			3374: dout = 12'h000;
			3375: dout = 12'h000;
			3376: dout = 12'h000;
			3377: dout = 12'ha61;
			3378: dout = 12'hf92;
			3379: dout = 12'hf82;
			3380: dout = 12'hc71;
			3381: dout = 12'h100;
			3382: dout = 12'h000;
			3383: dout = 12'h000;
			3384: dout = 12'h000;
			3385: dout = 12'h000;
			3386: dout = 12'h000;
			3387: dout = 12'h520;
			3388: dout = 12'h210;
			3389: dout = 12'h000;
			3390: dout = 12'h310;
			3391: dout = 12'h100;
			3392: dout = 12'h310;
			3393: dout = 12'h000;
			3394: dout = 12'h000;
			3395: dout = 12'h000;
			3396: dout = 12'h000;
			3397: dout = 12'h000;
			3398: dout = 12'h000;
			3399: dout = 12'h000;

			3400: dout = 12'h000;
			3401: dout = 12'h000;
			3402: dout = 12'h000;
			3403: dout = 12'h000;
			3404: dout = 12'h000;
			3405: dout = 12'h000;
			3406: dout = 12'h000;
			3407: dout = 12'h000;
			3408: dout = 12'h000;
			3409: dout = 12'h000;
			3410: dout = 12'h000;
			3411: dout = 12'h000;
			3412: dout = 12'h000;
			3413: dout = 12'h000;
			3414: dout = 12'h000;
			3415: dout = 12'h000;
			3416: dout = 12'h420;
			3417: dout = 12'h000;
			3418: dout = 12'hd62;
			3419: dout = 12'h631;
			3420: dout = 12'h100;
			3421: dout = 12'h000;
			3422: dout = 12'h000;
			3423: dout = 12'h000;
			3424: dout = 12'h000;
			3425: dout = 12'h000;
			3426: dout = 12'h000;
			3427: dout = 12'h000;
			3428: dout = 12'h000;
			3429: dout = 12'h000;
			3430: dout = 12'h000;
			3431: dout = 12'h000;
			3432: dout = 12'h000;
			3433: dout = 12'h520;
			3434: dout = 12'h100;
			3435: dout = 12'h000;
			3436: dout = 12'h000;
			3437: dout = 12'h000;
			3438: dout = 12'h000;
			3439: dout = 12'h000;

			3440: dout = 12'h000;
			3441: dout = 12'h000;
			3442: dout = 12'h000;
			3443: dout = 12'h000;
			3444: dout = 12'h000;
			3445: dout = 12'h000;
			3446: dout = 12'h000;
			3447: dout = 12'h000;
			3448: dout = 12'h000;
			3449: dout = 12'h000;
			3450: dout = 12'h000;
			3451: dout = 12'h000;
			3452: dout = 12'h000;
			3453: dout = 12'h000;
			3454: dout = 12'h000;
			3455: dout = 12'h000;
			3456: dout = 12'h310;
			3457: dout = 12'h000;
			3458: dout = 12'h310;
			3459: dout = 12'h000;
			3460: dout = 12'h000;
			3461: dout = 12'h000;
			3462: dout = 12'h000;
			3463: dout = 12'h000;
			3464: dout = 12'h000;
			3465: dout = 12'h000;
			3466: dout = 12'h000;
			3467: dout = 12'h000;
			3468: dout = 12'h000;
			3469: dout = 12'h000;
			3470: dout = 12'h000;
			3471: dout = 12'h000;
			3472: dout = 12'h000;
			3473: dout = 12'h000;
			3474: dout = 12'h000;
			3475: dout = 12'h000;
			3476: dout = 12'h000;
			3477: dout = 12'h000;
			3478: dout = 12'h000;
			3479: dout = 12'h000;

			3480: dout = 12'h000;
			3481: dout = 12'h000;
			3482: dout = 12'h000;
			3483: dout = 12'h000;
			3484: dout = 12'h000;
			3485: dout = 12'h000;
			3486: dout = 12'h000;
			3487: dout = 12'h000;
			3488: dout = 12'h000;
			3489: dout = 12'h000;
			3490: dout = 12'h000;
			3491: dout = 12'h000;
			3492: dout = 12'h000;
			3493: dout = 12'h000;
			3494: dout = 12'h000;
			3495: dout = 12'h000;
			3496: dout = 12'h000;
			3497: dout = 12'h000;
			3498: dout = 12'h000;
			3499: dout = 12'h000;
			3500: dout = 12'h000;
			3501: dout = 12'h000;
			3502: dout = 12'h000;
			3503: dout = 12'h000;
			3504: dout = 12'h000;
			3505: dout = 12'h000;
			3506: dout = 12'h000;
			3507: dout = 12'h000;
			3508: dout = 12'h000;
			3509: dout = 12'h000;
			3510: dout = 12'h000;
			3511: dout = 12'h000;
			3512: dout = 12'h000;
			3513: dout = 12'h000;
			3514: dout = 12'h000;
			3515: dout = 12'h000;
			3516: dout = 12'h000;
			3517: dout = 12'h000;
			3518: dout = 12'h000;
			3519: dout = 12'h000;

			3520: dout = 12'h000;
			3521: dout = 12'h000;
			3522: dout = 12'h000;
			3523: dout = 12'h000;
			3524: dout = 12'h000;
			3525: dout = 12'h114;
			3526: dout = 12'h44d;
			3527: dout = 12'h34c;
			3528: dout = 12'h34c;
			3529: dout = 12'h34c;
			3530: dout = 12'h34c;
			3531: dout = 12'h34c;
			3532: dout = 12'h34b;
			3533: dout = 12'h113;
			3534: dout = 12'h000;
			3535: dout = 12'h000;
			3536: dout = 12'h000;
			3537: dout = 12'h000;

			3538: dout = 12'h000;
			3539: dout = 12'h000;
			3540: dout = 12'h000;
			3541: dout = 12'h000;
			3542: dout = 12'h115;
			3543: dout = 12'h34a;
			3544: dout = 12'h47e;
			3545: dout = 12'h46d;
			3546: dout = 12'h46d;
			3547: dout = 12'h46d;
			3548: dout = 12'h46d;
			3549: dout = 12'h46d;
			3550: dout = 12'h46d;
			3551: dout = 12'h239;
			3552: dout = 12'h114;
			3553: dout = 12'h000;
			3554: dout = 12'h000;
			3555: dout = 12'h000;

			3556: dout = 12'h000;
			3557: dout = 12'h000;
			3558: dout = 12'h001;
			3559: dout = 12'h115;
			3560: dout = 12'h34b;
			3561: dout = 12'h46e;
			3562: dout = 12'h48e;
			3563: dout = 12'h48e;
			3564: dout = 12'h48e;
			3565: dout = 12'h48e;
			3566: dout = 12'h7ae;
			3567: dout = 12'h6ae;
			3568: dout = 12'h48e;
			3569: dout = 12'h46e;
			3570: dout = 12'h34a;
			3571: dout = 12'h113;
			3572: dout = 12'h001;
			3573: dout = 12'h000;

			3574: dout = 12'h000;
			3575: dout = 12'h001;
			3576: dout = 12'h126;
			3577: dout = 12'h45e;
			3578: dout = 12'h47e;
			3579: dout = 12'h48e;
			3580: dout = 12'h48e;
			3581: dout = 12'h48e;
			3582: dout = 12'h58e;
			3583: dout = 12'h69e;
			3584: dout = 12'hdef;
			3585: dout = 12'hbdf;
			3586: dout = 12'h48e;
			3587: dout = 12'h48e;
			3588: dout = 12'h47e;
			3589: dout = 12'h34c;
			3590: dout = 12'h114;
			3591: dout = 12'h001;

			3592: dout = 12'h001;
			3593: dout = 12'h228;
			3594: dout = 12'h35c;
			3595: dout = 12'h48e;
			3596: dout = 12'h48e;
			3597: dout = 12'h48e;
			3598: dout = 12'h48e;
			3599: dout = 12'h48e;
			3600: dout = 12'h8ae;
			3601: dout = 12'heff;
			3602: dout = 12'hfff;
			3603: dout = 12'hbdf;
			3604: dout = 12'h37e;
			3605: dout = 12'h48e;
			3606: dout = 12'h48e;
			3607: dout = 12'h47e;
			3608: dout = 12'h34c;
			3609: dout = 12'h226;

			3610: dout = 12'h001;
			3611: dout = 12'h33a;
			3612: dout = 12'h46d;
			3613: dout = 12'h48e;
			3614: dout = 12'h48e;
			3615: dout = 12'h48e;
			3616: dout = 12'h48e;
			3617: dout = 12'h48e;
			3618: dout = 12'h59e;
			3619: dout = 12'h7ae;
			3620: dout = 12'h7ae;
			3621: dout = 12'h9bf;
			3622: dout = 12'hbdf;
			3623: dout = 12'h69e;
			3624: dout = 12'h48e;
			3625: dout = 12'h48e;
			3626: dout = 12'h45d;
			3627: dout = 12'h227;

			3628: dout = 12'h001;
			3629: dout = 12'h339;
			3630: dout = 12'h45d;
			3631: dout = 12'h48e;
			3632: dout = 12'h48e;
			3633: dout = 12'h48e;
			3634: dout = 12'h48e;
			3635: dout = 12'h48e;
			3636: dout = 12'h48e;
			3637: dout = 12'h48e;
			3638: dout = 12'h48e;
			3639: dout = 12'h7ae;
			3640: dout = 12'hbdf;
			3641: dout = 12'h69e;
			3642: dout = 12'h48e;
			3643: dout = 12'h48e;
			3644: dout = 12'h45d;
			3645: dout = 12'h227;

			3646: dout = 12'h001;
			3647: dout = 12'h339;
			3648: dout = 12'h45d;
			3649: dout = 12'h48e;
			3650: dout = 12'h48e;
			3651: dout = 12'h48e;
			3652: dout = 12'h48e;
			3653: dout = 12'h48e;
			3654: dout = 12'h48e;
			3655: dout = 12'h48e;
			3656: dout = 12'h48e;
			3657: dout = 12'h48e;
			3658: dout = 12'h48e;
			3659: dout = 12'h48e;
			3660: dout = 12'h48e;
			3661: dout = 12'h48e;
			3662: dout = 12'h45d;
			3663: dout = 12'h227;

			3664: dout = 12'h001;
			3665: dout = 12'h339;
			3666: dout = 12'h45d;
			3667: dout = 12'h48e;
			3668: dout = 12'h48e;
			3669: dout = 12'h48e;
			3670: dout = 12'h48e;
			3671: dout = 12'h48e;
			3672: dout = 12'h48e;
			3673: dout = 12'h48e;
			3674: dout = 12'h48e;
			3675: dout = 12'h48e;
			3676: dout = 12'h48e;
			3677: dout = 12'h48e;
			3678: dout = 12'h48e;
			3679: dout = 12'h48e;
			3680: dout = 12'h45d;
			3681: dout = 12'h227;

			3682: dout = 12'h001;
			3683: dout = 12'h339;
			3684: dout = 12'h45d;
			3685: dout = 12'h48e;
			3686: dout = 12'h48e;
			3687: dout = 12'h48e;
			3688: dout = 12'h48e;
			3689: dout = 12'h48e;
			3690: dout = 12'h48e;
			3691: dout = 12'h48e;
			3692: dout = 12'h48e;
			3693: dout = 12'h48e;
			3694: dout = 12'h48e;
			3695: dout = 12'h48e;
			3696: dout = 12'h48e;
			3697: dout = 12'h48e;
			3698: dout = 12'h45d;
			3699: dout = 12'h227;

			3700: dout = 12'h001;
			3701: dout = 12'h339;
			3702: dout = 12'h45d;
			3703: dout = 12'h48e;
			3704: dout = 12'h48e;
			3705: dout = 12'h48e;
			3706: dout = 12'h48e;
			3707: dout = 12'h48e;
			3708: dout = 12'h48e;
			3709: dout = 12'h48e;
			3710: dout = 12'h48e;
			3711: dout = 12'h48e;
			3712: dout = 12'h48e;
			3713: dout = 12'h48e;
			3714: dout = 12'h48e;
			3715: dout = 12'h48e;
			3716: dout = 12'h45d;
			3717: dout = 12'h227;

			3718: dout = 12'h001;
			3719: dout = 12'h33a;
			3720: dout = 12'h46e;
			3721: dout = 12'h48e;
			3722: dout = 12'h48e;
			3723: dout = 12'h48e;
			3724: dout = 12'h48e;
			3725: dout = 12'h48e;
			3726: dout = 12'h48e;
			3727: dout = 12'h48e;
			3728: dout = 12'h48e;
			3729: dout = 12'h48e;
			3730: dout = 12'h48e;
			3731: dout = 12'h48e;
			3732: dout = 12'h48e;
			3733: dout = 12'h48e;
			3734: dout = 12'h45e;
			3735: dout = 12'h228;

			3736: dout = 12'h000;
			3737: dout = 12'h000;
			3738: dout = 12'h114;
			3739: dout = 12'h44d;
			3740: dout = 12'h47e;
			3741: dout = 12'h48e;
			3742: dout = 12'h48e;
			3743: dout = 12'h48e;
			3744: dout = 12'h48e;
			3745: dout = 12'h48e;
			3746: dout = 12'h48e;
			3747: dout = 12'h48e;
			3748: dout = 12'h48e;
			3749: dout = 12'h48e;
			3750: dout = 12'h46d;
			3751: dout = 12'h33b;
			3752: dout = 12'h002;
			3753: dout = 12'h000;

			3754: dout = 12'h000;
			3755: dout = 12'h000;
			3756: dout = 12'h002;
			3757: dout = 12'h226;
			3758: dout = 12'h35b;
			3759: dout = 12'h47e;
			3760: dout = 12'h48e;
			3761: dout = 12'h48e;
			3762: dout = 12'h48e;
			3763: dout = 12'h48e;
			3764: dout = 12'h48e;
			3765: dout = 12'h48e;
			3766: dout = 12'h48e;
			3767: dout = 12'h46e;
			3768: dout = 12'h34a;
			3769: dout = 12'h114;
			3770: dout = 12'h001;
			3771: dout = 12'h000;

			3772: dout = 12'h000;
			3773: dout = 12'h000;
			3774: dout = 12'h000;
			3775: dout = 12'h001;
			3776: dout = 12'h226;
			3777: dout = 12'h34a;
			3778: dout = 12'h47e;
			3779: dout = 12'h48e;
			3780: dout = 12'h48e;
			3781: dout = 12'h48e;
			3782: dout = 12'h48e;
			3783: dout = 12'h47e;
			3784: dout = 12'h46d;
			3785: dout = 12'h34a;
			3786: dout = 12'h115;
			3787: dout = 12'h000;
			3788: dout = 12'h000;
			3789: dout = 12'h000;

			3790: dout = 12'h000;
			3791: dout = 12'h000;
			3792: dout = 12'h000;
			3793: dout = 12'h000;
			3794: dout = 12'h000;
			3795: dout = 12'h113;
			3796: dout = 12'h34b;
			3797: dout = 12'h47d;
			3798: dout = 12'h48e;
			3799: dout = 12'h47e;
			3800: dout = 12'h48e;
			3801: dout = 12'h46d;
			3802: dout = 12'h33a;
			3803: dout = 12'h002;
			3804: dout = 12'h000;
			3805: dout = 12'h000;
			3806: dout = 12'h000;
			3807: dout = 12'h000;

			3808: dout = 12'h000;
			3809: dout = 12'h000;
			3810: dout = 12'h000;
			3811: dout = 12'h000;
			3812: dout = 12'h000;
			3813: dout = 12'h000;
			3814: dout = 12'h113;
			3815: dout = 12'h34b;
			3816: dout = 12'h45d;
			3817: dout = 12'h45d;
			3818: dout = 12'h45d;
			3819: dout = 12'h239;
			3820: dout = 12'h001;
			3821: dout = 12'h000;
			3822: dout = 12'h000;
			3823: dout = 12'h000;
			3824: dout = 12'h000;
			3825: dout = 12'h000;

			3826: dout = 12'h000;
			3827: dout = 12'h000;
			3828: dout = 12'h000;
			3829: dout = 12'h000;
			3830: dout = 12'h000;
			3831: dout = 12'h000;
			3832: dout = 12'h000;
			3833: dout = 12'h002;
			3834: dout = 12'h227;
			3835: dout = 12'h34c;
			3836: dout = 12'h125;
			3837: dout = 12'h002;
			3838: dout = 12'h000;
			3839: dout = 12'h000;
			3840: dout = 12'h000;
			3841: dout = 12'h000;
			3842: dout = 12'h000;
			3843: dout = 12'h000;

			3844: dout = 12'h000;
			3845: dout = 12'h000;
			3846: dout = 12'h000;
			3847: dout = 12'h000;
			3848: dout = 12'h000;
			3849: dout = 12'h000;
			3850: dout = 12'h000;
			3851: dout = 12'h000;
			3852: dout = 12'h114;
			3853: dout = 12'h34c;
			3854: dout = 12'h113;
			3855: dout = 12'h000;
			3856: dout = 12'h000;
			3857: dout = 12'h000;
			3858: dout = 12'h000;
			3859: dout = 12'h000;
			3860: dout = 12'h000;
			3861: dout = 12'h000;

			3862: dout = 12'h000;
			3863: dout = 12'h000;
			3864: dout = 12'h000;
			3865: dout = 12'h000;
			3866: dout = 12'h000;
			3867: dout = 12'h000;
			3868: dout = 12'h001;
			3869: dout = 12'h001;
			3870: dout = 12'h115;
			3871: dout = 12'h33a;
			3872: dout = 12'h012;
			3873: dout = 12'h000;
			3874: dout = 12'h000;
			3875: dout = 12'h000;
			3876: dout = 12'h000;
			3877: dout = 12'h000;
			3878: dout = 12'h000;
			3879: dout = 12'h000;

			3880: dout = 12'h000;
			3881: dout = 12'h000;
			3882: dout = 12'h000;
			3883: dout = 12'h000;
			3884: dout = 12'h000;
			3885: dout = 12'h114;
			3886: dout = 12'h34c;
			3887: dout = 12'h34c;
			3888: dout = 12'h228;
			3889: dout = 12'h002;
			3890: dout = 12'h000;
			3891: dout = 12'h000;
			3892: dout = 12'h000;
			3893: dout = 12'h000;
			3894: dout = 12'h000;
			3895: dout = 12'h000;
			3896: dout = 12'h000;
			3897: dout = 12'h000;

			3898: dout = 12'h000;
			3899: dout = 12'h000;
			3900: dout = 12'h000;
			3901: dout = 12'h001;
			3902: dout = 12'h227;
			3903: dout = 12'h227;
			3904: dout = 12'h114;
			3905: dout = 12'h114;
			3906: dout = 12'h002;
			3907: dout = 12'h000;
			3908: dout = 12'h000;
			3909: dout = 12'h000;
			3910: dout = 12'h000;
			3911: dout = 12'h000;
			3912: dout = 12'h000;
			3913: dout = 12'h000;
			3914: dout = 12'h000;
			3915: dout = 12'h000;

			3916: dout = 12'h000;
			3917: dout = 12'h000;
			3918: dout = 12'h002;
			3919: dout = 12'h126;
			3920: dout = 12'h227;
			3921: dout = 12'h115;
			3922: dout = 12'h000;
			3923: dout = 12'h000;
			3924: dout = 12'h000;
			3925: dout = 12'h000;
			3926: dout = 12'h000;
			3927: dout = 12'h000;
			3928: dout = 12'h000;
			3929: dout = 12'h000;
			3930: dout = 12'h000;
			3931: dout = 12'h000;
			3932: dout = 12'h000;
			3933: dout = 12'h000;

			3934: dout = 12'h000;
			3935: dout = 12'h000;
			3936: dout = 12'h114;
			3937: dout = 12'h34c;
			3938: dout = 12'h113;
			3939: dout = 12'h000;
			3940: dout = 12'h000;
			3941: dout = 12'h000;
			3942: dout = 12'h000;
			3943: dout = 12'h000;
			3944: dout = 12'h000;
			3945: dout = 12'h000;
			3946: dout = 12'h000;
			3947: dout = 12'h000;
			3948: dout = 12'h000;
			3949: dout = 12'h000;
			3950: dout = 12'h000;
			3951: dout = 12'h000;

			3952: dout = 12'h000;
			3953: dout = 12'h000;
			3954: dout = 12'h000;
			3955: dout = 12'h000;
			3956: dout = 12'h000;
			3957: dout = 12'h001;
			3958: dout = 12'h113;
			3959: dout = 12'h113;
			3960: dout = 12'h113;
			3961: dout = 12'h113;
			3962: dout = 12'h113;
			3963: dout = 12'h113;
			3964: dout = 12'h013;
			3965: dout = 12'h001;
			3966: dout = 12'h000;
			3967: dout = 12'h000;
			3968: dout = 12'h000;
			3969: dout = 12'h000;

			3970: dout = 12'h000;
			3971: dout = 12'h000;
			3972: dout = 12'h000;
			3973: dout = 12'h000;
			3974: dout = 12'h115;
			3975: dout = 12'h34a;
			3976: dout = 12'h47e;
			3977: dout = 12'h46d;
			3978: dout = 12'h46d;
			3979: dout = 12'h46d;
			3980: dout = 12'h46d;
			3981: dout = 12'h46d;
			3982: dout = 12'h46d;
			3983: dout = 12'h239;
			3984: dout = 12'h114;
			3985: dout = 12'h000;
			3986: dout = 12'h000;
			3987: dout = 12'h000;

			3988: dout = 12'h000;
			3989: dout = 12'h000;
			3990: dout = 12'h001;
			3991: dout = 12'h115;
			3992: dout = 12'h34b;
			3993: dout = 12'h46e;
			3994: dout = 12'h48e;
			3995: dout = 12'h48e;
			3996: dout = 12'h48e;
			3997: dout = 12'h48e;
			3998: dout = 12'h7ae;
			3999: dout = 12'h6ae;
			4000: dout = 12'h48e;
			4001: dout = 12'h46e;
			4002: dout = 12'h34a;
			4003: dout = 12'h013;
			4004: dout = 12'h000;
			4005: dout = 12'h000;

			4006: dout = 12'h000;
			4007: dout = 12'h001;
			4008: dout = 12'h126;
			4009: dout = 12'h45e;
			4010: dout = 12'h47e;
			4011: dout = 12'h48e;
			4012: dout = 12'h48e;
			4013: dout = 12'h48e;
			4014: dout = 12'h58e;
			4015: dout = 12'h69e;
			4016: dout = 12'hdef;
			4017: dout = 12'hbdf;
			4018: dout = 12'h48e;
			4019: dout = 12'h48e;
			4020: dout = 12'h47e;
			4021: dout = 12'h34b;
			4022: dout = 12'h001;
			4023: dout = 12'h000;

			4024: dout = 12'h000;
			4025: dout = 12'h115;
			4026: dout = 12'h35c;
			4027: dout = 12'h48e;
			4028: dout = 12'h48e;
			4029: dout = 12'h48e;
			4030: dout = 12'h48e;
			4031: dout = 12'h48e;
			4032: dout = 12'h8ae;
			4033: dout = 12'heff;
			4034: dout = 12'hfff;
			4035: dout = 12'hbdf;
			4036: dout = 12'h37e;
			4037: dout = 12'h48e;
			4038: dout = 12'h48e;
			4039: dout = 12'h47e;
			4040: dout = 12'h226;
			4041: dout = 12'h000;

			4042: dout = 12'h000;
			4043: dout = 12'h226;
			4044: dout = 12'h46d;
			4045: dout = 12'h48e;
			4046: dout = 12'h48e;
			4047: dout = 12'h48e;
			4048: dout = 12'h48e;
			4049: dout = 12'h48e;
			4050: dout = 12'h59e;
			4051: dout = 12'h7ae;
			4052: dout = 12'h7ae;
			4053: dout = 12'h9bf;
			4054: dout = 12'hbdf;
			4055: dout = 12'h69e;
			4056: dout = 12'h48e;
			4057: dout = 12'h48e;
			4058: dout = 12'h236;
			4059: dout = 12'h000;

			4060: dout = 12'h000;
			4061: dout = 12'h226;
			4062: dout = 12'h45d;
			4063: dout = 12'h48e;
			4064: dout = 12'h48e;
			4065: dout = 12'h48e;
			4066: dout = 12'h48e;
			4067: dout = 12'h48e;
			4068: dout = 12'h48e;
			4069: dout = 12'h48e;
			4070: dout = 12'h48e;
			4071: dout = 12'h7ae;
			4072: dout = 12'hbdf;
			4073: dout = 12'h69e;
			4074: dout = 12'h48e;
			4075: dout = 12'h48e;
			4076: dout = 12'h236;
			4077: dout = 12'h000;

			4078: dout = 12'h000;
			4079: dout = 12'h226;
			4080: dout = 12'h45d;
			4081: dout = 12'h48e;
			4082: dout = 12'h48e;
			4083: dout = 12'h48e;
			4084: dout = 12'h48e;
			4085: dout = 12'h48e;
			4086: dout = 12'h48e;
			4087: dout = 12'h48e;
			4088: dout = 12'h48e;
			4089: dout = 12'h48e;
			4090: dout = 12'h48e;
			4091: dout = 12'h48e;
			4092: dout = 12'h48e;
			4093: dout = 12'h48e;
			4094: dout = 12'h236;
			4095: dout = 12'h000;

			4096: dout = 12'h000;
			4097: dout = 12'h226;
			4098: dout = 12'h45d;
			4099: dout = 12'h48e;
			4100: dout = 12'h48e;
			4101: dout = 12'h48e;
			4102: dout = 12'h48e;
			4103: dout = 12'h48e;
			4104: dout = 12'h48e;
			4105: dout = 12'h48e;
			4106: dout = 12'h48e;
			4107: dout = 12'h48e;
			4108: dout = 12'h48e;
			4109: dout = 12'h48e;
			4110: dout = 12'h48e;
			4111: dout = 12'h48e;
			4112: dout = 12'h236;
			4113: dout = 12'h000;

			4114: dout = 12'h000;
			4115: dout = 12'h226;
			4116: dout = 12'h45d;
			4117: dout = 12'h48e;
			4118: dout = 12'h48e;
			4119: dout = 12'h48e;
			4120: dout = 12'h48e;
			4121: dout = 12'h48e;
			4122: dout = 12'h48e;
			4123: dout = 12'h48e;
			4124: dout = 12'h48e;
			4125: dout = 12'h48e;
			4126: dout = 12'h48e;
			4127: dout = 12'h48e;
			4128: dout = 12'h48e;
			4129: dout = 12'h48e;
			4130: dout = 12'h236;
			4131: dout = 12'h000;

			4132: dout = 12'h000;
			4133: dout = 12'h226;
			4134: dout = 12'h45d;
			4135: dout = 12'h48e;
			4136: dout = 12'h48e;
			4137: dout = 12'h48e;
			4138: dout = 12'h48e;
			4139: dout = 12'h48e;
			4140: dout = 12'h48e;
			4141: dout = 12'h48e;
			4142: dout = 12'h48e;
			4143: dout = 12'h48e;
			4144: dout = 12'h48e;
			4145: dout = 12'h48e;
			4146: dout = 12'h48e;
			4147: dout = 12'h48e;
			4148: dout = 12'h236;
			4149: dout = 12'h000;

			4150: dout = 12'h000;
			4151: dout = 12'h227;
			4152: dout = 12'h46e;
			4153: dout = 12'h48e;
			4154: dout = 12'h48e;
			4155: dout = 12'h48e;
			4156: dout = 12'h48e;
			4157: dout = 12'h48e;
			4158: dout = 12'h48e;
			4159: dout = 12'h48e;
			4160: dout = 12'h48e;
			4161: dout = 12'h48e;
			4162: dout = 12'h48e;
			4163: dout = 12'h48e;
			4164: dout = 12'h48e;
			4165: dout = 12'h48e;
			4166: dout = 12'h237;
			4167: dout = 12'h000;

			4168: dout = 12'h000;
			4169: dout = 12'h000;
			4170: dout = 12'h113;
			4171: dout = 12'h44d;
			4172: dout = 12'h47e;
			4173: dout = 12'h48e;
			4174: dout = 12'h48e;
			4175: dout = 12'h48e;
			4176: dout = 12'h48e;
			4177: dout = 12'h48e;
			4178: dout = 12'h48e;
			4179: dout = 12'h48e;
			4180: dout = 12'h48e;
			4181: dout = 12'h48e;
			4182: dout = 12'h46d;
			4183: dout = 12'h33a;
			4184: dout = 12'h002;
			4185: dout = 12'h000;

			4186: dout = 12'h000;
			4187: dout = 12'h000;
			4188: dout = 12'h000;
			4189: dout = 12'h226;
			4190: dout = 12'h35b;
			4191: dout = 12'h47e;
			4192: dout = 12'h48e;
			4193: dout = 12'h48e;
			4194: dout = 12'h48e;
			4195: dout = 12'h48e;
			4196: dout = 12'h48e;
			4197: dout = 12'h48e;
			4198: dout = 12'h48e;
			4199: dout = 12'h46e;
			4200: dout = 12'h34a;
			4201: dout = 12'h114;
			4202: dout = 12'h000;
			4203: dout = 12'h000;

			4204: dout = 12'h000;
			4205: dout = 12'h000;
			4206: dout = 12'h000;
			4207: dout = 12'h001;
			4208: dout = 12'h226;
			4209: dout = 12'h34a;
			4210: dout = 12'h47e;
			4211: dout = 12'h48e;
			4212: dout = 12'h48e;
			4213: dout = 12'h48e;
			4214: dout = 12'h48e;
			4215: dout = 12'h47e;
			4216: dout = 12'h46d;
			4217: dout = 12'h34a;
			4218: dout = 12'h115;
			4219: dout = 12'h000;
			4220: dout = 12'h000;
			4221: dout = 12'h000;

			4222: dout = 12'h000;
			4223: dout = 12'h000;
			4224: dout = 12'h000;
			4225: dout = 12'h000;
			4226: dout = 12'h000;
			4227: dout = 12'h113;
			4228: dout = 12'h34b;
			4229: dout = 12'h47d;
			4230: dout = 12'h48e;
			4231: dout = 12'h47e;
			4232: dout = 12'h48e;
			4233: dout = 12'h46d;
			4234: dout = 12'h33a;
			4235: dout = 12'h002;
			4236: dout = 12'h000;
			4237: dout = 12'h000;
			4238: dout = 12'h000;
			4239: dout = 12'h000;

			4240: dout = 12'h000;
			4241: dout = 12'h000;
			4242: dout = 12'h000;
			4243: dout = 12'h000;
			4244: dout = 12'h000;
			4245: dout = 12'h000;
			4246: dout = 12'h113;
			4247: dout = 12'h34b;
			4248: dout = 12'h45d;
			4249: dout = 12'h45d;
			4250: dout = 12'h45d;
			4251: dout = 12'h239;
			4252: dout = 12'h001;
			4253: dout = 12'h000;
			4254: dout = 12'h000;
			4255: dout = 12'h000;
			4256: dout = 12'h000;
			4257: dout = 12'h000;

			4258: dout = 12'h000;
			4259: dout = 12'h000;
			4260: dout = 12'h000;
			4261: dout = 12'h000;
			4262: dout = 12'h000;
			4263: dout = 12'h000;
			4264: dout = 12'h000;
			4265: dout = 12'h002;
			4266: dout = 12'h227;
			4267: dout = 12'h34c;
			4268: dout = 12'h125;
			4269: dout = 12'h002;
			4270: dout = 12'h000;
			4271: dout = 12'h000;
			4272: dout = 12'h000;
			4273: dout = 12'h000;
			4274: dout = 12'h000;
			4275: dout = 12'h000;

			4276: dout = 12'h000;
			4277: dout = 12'h000;
			4278: dout = 12'h000;
			4279: dout = 12'h000;
			4280: dout = 12'h000;
			4281: dout = 12'h000;
			4282: dout = 12'h000;
			4283: dout = 12'h000;
			4284: dout = 12'h114;
			4285: dout = 12'h34c;
			4286: dout = 12'h113;
			4287: dout = 12'h000;
			4288: dout = 12'h000;
			4289: dout = 12'h000;
			4290: dout = 12'h000;
			4291: dout = 12'h000;
			4292: dout = 12'h000;
			4293: dout = 12'h000;

			4294: dout = 12'h000;
			4295: dout = 12'h000;
			4296: dout = 12'h000;
			4297: dout = 12'h000;
			4298: dout = 12'h000;
			4299: dout = 12'h000;
			4300: dout = 12'h000;
			4301: dout = 12'h113;
			4302: dout = 12'h239;
			4303: dout = 12'h33a;
			4304: dout = 12'h012;
			4305: dout = 12'h000;
			4306: dout = 12'h000;
			4307: dout = 12'h000;
			4308: dout = 12'h000;
			4309: dout = 12'h000;
			4310: dout = 12'h000;
			4311: dout = 12'h000;

			4312: dout = 12'h000;
			4313: dout = 12'h000;
			4314: dout = 12'h000;
			4315: dout = 12'h000;
			4316: dout = 12'h000;
			4317: dout = 12'h000;
			4318: dout = 12'h000;
			4319: dout = 12'h228;
			4320: dout = 12'h33a;
			4321: dout = 12'h002;
			4322: dout = 12'h000;
			4323: dout = 12'h000;
			4324: dout = 12'h000;
			4325: dout = 12'h000;
			4326: dout = 12'h000;
			4327: dout = 12'h000;
			4328: dout = 12'h000;
			4329: dout = 12'h000;

			4330: dout = 12'h000;
			4331: dout = 12'h000;
			4332: dout = 12'h000;
			4333: dout = 12'h000;
			4334: dout = 12'h000;
			4335: dout = 12'h000;
			4336: dout = 12'h126;
			4337: dout = 12'h226;
			4338: dout = 12'h002;
			4339: dout = 12'h000;
			4340: dout = 12'h000;
			4341: dout = 12'h000;
			4342: dout = 12'h000;
			4343: dout = 12'h000;
			4344: dout = 12'h000;
			4345: dout = 12'h000;
			4346: dout = 12'h000;
			4347: dout = 12'h000;

			4348: dout = 12'h000;
			4349: dout = 12'h000;
			4350: dout = 12'h000;
			4351: dout = 12'h000;
			4352: dout = 12'h000;
			4353: dout = 12'h114;
			4354: dout = 12'h114;
			4355: dout = 12'h000;
			4356: dout = 12'h000;
			4357: dout = 12'h000;
			4358: dout = 12'h000;
			4359: dout = 12'h000;
			4360: dout = 12'h000;
			4361: dout = 12'h000;
			4362: dout = 12'h000;
			4363: dout = 12'h000;
			4364: dout = 12'h000;
			4365: dout = 12'h000;

			4366: dout = 12'h000;
			4367: dout = 12'h000;
			4368: dout = 12'h000;
			4369: dout = 12'h000;
			4370: dout = 12'h000;
			4371: dout = 12'h002;
			4372: dout = 12'h000;
			4373: dout = 12'h000;
			4374: dout = 12'h000;
			4375: dout = 12'h000;
			4376: dout = 12'h000;
			4377: dout = 12'h000;
			4378: dout = 12'h000;
			4379: dout = 12'h000;
			4380: dout = 12'h000;
			4381: dout = 12'h000;
			4382: dout = 12'h000;
			4383: dout = 12'h000;

			4384: dout = 12'h000;
			4385: dout = 12'h812;
			4386: dout = 12'he33;
			4387: dout = 12'hd33;
			4388: dout = 12'hd33;
			4389: dout = 12'hd33;
			4390: dout = 12'ha23;
			4391: dout = 12'h000;

			4392: dout = 12'h803;
			4393: dout = 12'hfa2;
			4394: dout = 12'hfe1;
			4395: dout = 12'hfe1;
			4396: dout = 12'hfe1;
			4397: dout = 12'hfe1;
			4398: dout = 12'hfc2;
			4399: dout = 12'hb24;

			4400: dout = 12'h000;
			4401: dout = 12'h712;
			4402: dout = 12'hd33;
			4403: dout = 12'hc23;
			4404: dout = 12'hc23;
			4405: dout = 12'hd33;
			4406: dout = 12'h913;
			4407: dout = 12'h000;

			4408: dout = 12'h000;
			4409: dout = 12'h000;
			4410: dout = 12'h000;
			4411: dout = 12'h000;
			4412: dout = 12'h000;
			4413: dout = 12'h000;
			4414: dout = 12'h000;
			4415: dout = 12'h000;
			4416: dout = 12'h000;
			4417: dout = 12'h000;
			4418: dout = 12'h000;
			4419: dout = 12'h000;
			4420: dout = 12'h000;
			4421: dout = 12'h000;
			4422: dout = 12'h000;
			4423: dout = 12'h000;
			4424: dout = 12'h000;
			4425: dout = 12'h000;
			4426: dout = 12'h000;
			4427: dout = 12'h000;
			4428: dout = 12'h000;
			4429: dout = 12'h000;
			4430: dout = 12'h000;
			4431: dout = 12'h000;
			4432: dout = 12'h000;
			4433: dout = 12'h000;
			4434: dout = 12'h000;
			4435: dout = 12'h000;
			4436: dout = 12'h000;
			4437: dout = 12'h000;
			4438: dout = 12'h000;
			4439: dout = 12'h000;
			4440: dout = 12'h000;
			4441: dout = 12'h000;
			4442: dout = 12'h000;
			4443: dout = 12'h000;
			4444: dout = 12'h000;
			4445: dout = 12'h000;
			4446: dout = 12'h000;
			4447: dout = 12'h000;
			4448: dout = 12'h000;
			4449: dout = 12'h000;
			4450: dout = 12'h000;
			4451: dout = 12'h000;
			4452: dout = 12'h000;
			4453: dout = 12'h000;
			4454: dout = 12'h000;
			4455: dout = 12'h000;
			4456: dout = 12'h000;
			4457: dout = 12'h000;
			4458: dout = 12'h000;
			4459: dout = 12'h000;
			4460: dout = 12'h000;
			4461: dout = 12'h000;
			4462: dout = 12'h000;
			4463: dout = 12'h000;
			4464: dout = 12'h000;
			4465: dout = 12'h000;
			4466: dout = 12'h000;
			4467: dout = 12'h000;
			4468: dout = 12'h000;
			4469: dout = 12'h000;
			4470: dout = 12'h000;
			4471: dout = 12'h000;
			4472: dout = 12'h000;
			4473: dout = 12'h000;
			4474: dout = 12'h000;
			4475: dout = 12'h000;
			4476: dout = 12'h000;
			4477: dout = 12'h000;
			4478: dout = 12'h000;
			4479: dout = 12'h000;
			4480: dout = 12'h000;
			4481: dout = 12'h000;
			4482: dout = 12'h000;
			4483: dout = 12'h000;
			4484: dout = 12'h000;
			4485: dout = 12'h000;
			4486: dout = 12'h000;
			4487: dout = 12'h000;
			4488: dout = 12'h000;
			4489: dout = 12'h000;
			4490: dout = 12'h000;
			4491: dout = 12'h000;
			4492: dout = 12'h000;
			4493: dout = 12'h000;
			4494: dout = 12'h000;
			4495: dout = 12'h000;
			4496: dout = 12'h000;
			4497: dout = 12'h000;
			4498: dout = 12'h000;
			4499: dout = 12'h000;
			4500: dout = 12'h000;
			4501: dout = 12'h000;
			4502: dout = 12'h000;
			4503: dout = 12'h000;
			4504: dout = 12'h000;
			4505: dout = 12'h000;
			4506: dout = 12'h000;
			4507: dout = 12'h000;
			4508: dout = 12'h000;
			4509: dout = 12'h000;
			4510: dout = 12'h000;
			4511: dout = 12'h000;
			4512: dout = 12'h000;
			4513: dout = 12'h000;
			4514: dout = 12'h000;
			4515: dout = 12'h000;
			4516: dout = 12'h000;
			4517: dout = 12'h000;
			4518: dout = 12'h000;
			4519: dout = 12'h000;
			4520: dout = 12'h000;
			4521: dout = 12'h000;
			4522: dout = 12'h000;
			4523: dout = 12'h000;
			4524: dout = 12'h000;
			4525: dout = 12'h000;
			4526: dout = 12'h000;
			4527: dout = 12'h000;
			4528: dout = 12'h000;
			4529: dout = 12'h000;
			4530: dout = 12'h000;
			4531: dout = 12'h000;
			4532: dout = 12'h000;
			4533: dout = 12'h000;
			4534: dout = 12'h000;
			4535: dout = 12'h000;
			4536: dout = 12'h000;
			4537: dout = 12'h000;
			4538: dout = 12'h000;
			4539: dout = 12'h000;
			4540: dout = 12'h000;
			4541: dout = 12'h000;
			4542: dout = 12'h000;
			4543: dout = 12'h000;
			4544: dout = 12'h000;
			4545: dout = 12'h000;
			4546: dout = 12'h000;
			4547: dout = 12'h000;
			4548: dout = 12'h000;
			4549: dout = 12'h000;
			4550: dout = 12'h000;
			4551: dout = 12'h000;
			4552: dout = 12'h000;
			4553: dout = 12'h000;
			4554: dout = 12'h000;
			4555: dout = 12'h000;
			4556: dout = 12'h000;
			4557: dout = 12'h000;

			4558: dout = 12'h000;
			4559: dout = 12'h000;
			4560: dout = 12'h000;
			4561: dout = 12'h000;
			4562: dout = 12'h000;
			4563: dout = 12'h000;
			4564: dout = 12'h000;
			4565: dout = 12'h000;
			4566: dout = 12'h000;
			4567: dout = 12'h000;
			4568: dout = 12'h000;
			4569: dout = 12'h000;
			4570: dout = 12'h000;
			4571: dout = 12'h000;
			4572: dout = 12'h000;
			4573: dout = 12'h000;
			4574: dout = 12'h000;
			4575: dout = 12'h000;
			4576: dout = 12'h000;
			4577: dout = 12'h000;
			4578: dout = 12'h000;
			4579: dout = 12'h000;
			4580: dout = 12'h000;
			4581: dout = 12'h000;
			4582: dout = 12'h000;
			4583: dout = 12'h000;
			4584: dout = 12'h000;
			4585: dout = 12'h000;
			4586: dout = 12'h000;
			4587: dout = 12'h000;
			4588: dout = 12'h000;
			4589: dout = 12'h000;
			4590: dout = 12'h000;
			4591: dout = 12'h000;
			4592: dout = 12'h000;
			4593: dout = 12'h000;
			4594: dout = 12'h000;
			4595: dout = 12'h000;
			4596: dout = 12'h000;
			4597: dout = 12'h000;
			4598: dout = 12'h000;
			4599: dout = 12'h000;
			4600: dout = 12'h000;
			4601: dout = 12'h000;
			4602: dout = 12'h000;
			4603: dout = 12'h000;
			4604: dout = 12'h000;
			4605: dout = 12'h000;
			4606: dout = 12'h000;
			4607: dout = 12'h000;
			4608: dout = 12'h000;
			4609: dout = 12'h000;
			4610: dout = 12'h000;
			4611: dout = 12'h000;
			4612: dout = 12'h000;
			4613: dout = 12'h000;
			4614: dout = 12'h000;
			4615: dout = 12'h000;
			4616: dout = 12'h000;
			4617: dout = 12'h000;
			4618: dout = 12'h000;
			4619: dout = 12'h000;
			4620: dout = 12'h000;
			4621: dout = 12'h000;
			4622: dout = 12'h000;
			4623: dout = 12'h000;
			4624: dout = 12'h000;
			4625: dout = 12'h000;
			4626: dout = 12'h000;
			4627: dout = 12'h000;
			4628: dout = 12'h000;
			4629: dout = 12'h000;
			4630: dout = 12'h000;
			4631: dout = 12'h000;
			4632: dout = 12'h000;
			4633: dout = 12'h000;
			4634: dout = 12'h000;
			4635: dout = 12'h000;
			4636: dout = 12'h000;
			4637: dout = 12'h000;
			4638: dout = 12'h000;
			4639: dout = 12'h000;
			4640: dout = 12'h000;
			4641: dout = 12'h000;
			4642: dout = 12'h000;
			4643: dout = 12'h000;
			4644: dout = 12'h000;
			4645: dout = 12'h000;
			4646: dout = 12'h000;
			4647: dout = 12'h000;
			4648: dout = 12'h000;
			4649: dout = 12'h000;
			4650: dout = 12'h000;
			4651: dout = 12'h000;
			4652: dout = 12'h000;
			4653: dout = 12'h000;
			4654: dout = 12'h000;
			4655: dout = 12'h000;
			4656: dout = 12'h000;
			4657: dout = 12'h000;
			4658: dout = 12'h000;
			4659: dout = 12'h000;
			4660: dout = 12'h000;
			4661: dout = 12'h000;
			4662: dout = 12'h000;
			4663: dout = 12'h000;
			4664: dout = 12'h000;
			4665: dout = 12'h000;
			4666: dout = 12'h000;
			4667: dout = 12'h000;
			4668: dout = 12'h000;
			4669: dout = 12'h000;
			4670: dout = 12'h000;
			4671: dout = 12'h000;
			4672: dout = 12'h000;
			4673: dout = 12'h000;
			4674: dout = 12'h000;
			4675: dout = 12'h000;
			4676: dout = 12'h000;
			4677: dout = 12'h000;
			4678: dout = 12'h000;
			4679: dout = 12'h000;
			4680: dout = 12'h000;
			4681: dout = 12'h000;
			4682: dout = 12'h000;
			4683: dout = 12'h000;
			4684: dout = 12'h000;
			4685: dout = 12'h000;
			4686: dout = 12'h000;
			4687: dout = 12'h000;
			4688: dout = 12'h000;
			4689: dout = 12'h000;
			4690: dout = 12'h000;
			4691: dout = 12'h000;
			4692: dout = 12'h000;
			4693: dout = 12'h000;
			4694: dout = 12'h000;
			4695: dout = 12'h000;
			4696: dout = 12'h000;
			4697: dout = 12'h000;
			4698: dout = 12'h000;
			4699: dout = 12'h000;
			4700: dout = 12'h000;
			4701: dout = 12'h000;
			4702: dout = 12'h000;
			4703: dout = 12'h000;
			4704: dout = 12'h000;
			4705: dout = 12'h000;
			4706: dout = 12'h000;
			4707: dout = 12'h000;

			4708: dout = 12'h000;
			4709: dout = 12'h000;
			4710: dout = 12'h000;
			4711: dout = 12'h000;
			4712: dout = 12'h000;
			4713: dout = 12'h800;
			4714: dout = 12'hd00;
			4715: dout = 12'hc00;
			4716: dout = 12'hc00;
			4717: dout = 12'hc00;
			4718: dout = 12'hc00;
			4719: dout = 12'hc00;
			4720: dout = 12'hc00;
			4721: dout = 12'hc00;
			4722: dout = 12'hc00;
			4723: dout = 12'hc00;
			4724: dout = 12'hc00;
			4725: dout = 12'hc00;
			4726: dout = 12'hc00;
			4727: dout = 12'h200;
			4728: dout = 12'h000;
			4729: dout = 12'h000;
			4730: dout = 12'h000;
			4731: dout = 12'h500;
			4732: dout = 12'hd00;
			4733: dout = 12'hc00;
			4734: dout = 12'hc00;
			4735: dout = 12'hc00;
			4736: dout = 12'hc00;
			4737: dout = 12'hc00;
			4738: dout = 12'hd00;
			4739: dout = 12'h300;
			4740: dout = 12'h000;
			4741: dout = 12'h000;
			4742: dout = 12'h000;
			4743: dout = 12'h400;
			4744: dout = 12'hd00;
			4745: dout = 12'hc00;
			4746: dout = 12'ha00;
			4747: dout = 12'h000;
			4748: dout = 12'h000;
			4749: dout = 12'h000;
			4750: dout = 12'h000;
			4751: dout = 12'h000;
			4752: dout = 12'h000;
			4753: dout = 12'h000;
			4754: dout = 12'h000;
			4755: dout = 12'h300;
			4756: dout = 12'hd00;
			4757: dout = 12'hc00;
			4758: dout = 12'hc10;
			4759: dout = 12'h000;
			4760: dout = 12'h900;
			4761: dout = 12'hc00;
			4762: dout = 12'hc00;
			4763: dout = 12'hc00;
			4764: dout = 12'hc00;
			4765: dout = 12'hc00;
			4766: dout = 12'hc00;
			4767: dout = 12'hc00;
			4768: dout = 12'hc00;
			4769: dout = 12'hc00;
			4770: dout = 12'hc00;
			4771: dout = 12'hc00;
			4772: dout = 12'hc00;
			4773: dout = 12'hc00;
			4774: dout = 12'hd00;
			4775: dout = 12'h700;
			4776: dout = 12'h000;
			4777: dout = 12'h000;
			4778: dout = 12'h000;
			4779: dout = 12'h000;
			4780: dout = 12'h000;
			4781: dout = 12'h000;
			4782: dout = 12'h000;
			4783: dout = 12'h000;
			4784: dout = 12'h000;
			4785: dout = 12'h000;
			4786: dout = 12'h000;
			4787: dout = 12'h600;
			4788: dout = 12'hd00;
			4789: dout = 12'hc00;
			4790: dout = 12'hc00;
			4791: dout = 12'hc00;
			4792: dout = 12'hc00;
			4793: dout = 12'hc00;
			4794: dout = 12'hc00;
			4795: dout = 12'hc00;
			4796: dout = 12'hc00;
			4797: dout = 12'hc00;
			4798: dout = 12'hc00;
			4799: dout = 12'ha00;
			4800: dout = 12'h000;
			4801: dout = 12'h000;
			4802: dout = 12'h000;
			4803: dout = 12'h000;
			4804: dout = 12'hb10;
			4805: dout = 12'hc00;
			4806: dout = 12'hd00;
			4807: dout = 12'h300;
			4808: dout = 12'h000;
			4809: dout = 12'h000;
			4810: dout = 12'h000;
			4811: dout = 12'h000;
			4812: dout = 12'h000;
			4813: dout = 12'h000;
			4814: dout = 12'h000;
			4815: dout = 12'h000;
			4816: dout = 12'ha00;
			4817: dout = 12'hc00;
			4818: dout = 12'hd00;
			4819: dout = 12'h400;
			4820: dout = 12'h200;
			4821: dout = 12'hd00;
			4822: dout = 12'hc00;
			4823: dout = 12'hc00;
			4824: dout = 12'hc00;
			4825: dout = 12'hc00;
			4826: dout = 12'hc00;
			4827: dout = 12'hc00;
			4828: dout = 12'hc00;
			4829: dout = 12'hc00;
			4830: dout = 12'hc00;
			4831: dout = 12'hc00;
			4832: dout = 12'hc00;
			4833: dout = 12'hc00;
			4834: dout = 12'hc00;
			4835: dout = 12'hc00;
			4836: dout = 12'h000;
			4837: dout = 12'h800;
			4838: dout = 12'hd00;
			4839: dout = 12'hc00;
			4840: dout = 12'hc00;
			4841: dout = 12'hc00;
			4842: dout = 12'hc00;
			4843: dout = 12'hc00;
			4844: dout = 12'hc00;
			4845: dout = 12'hc00;
			4846: dout = 12'hc00;
			4847: dout = 12'hc00;
			4848: dout = 12'hc00;
			4849: dout = 12'hc00;
			4850: dout = 12'hc00;
			4851: dout = 12'h200;
			4852: dout = 12'h000;
			4853: dout = 12'h000;
			4854: dout = 12'h000;
			4855: dout = 12'h000;
			4856: dout = 12'h000;
			4857: dout = 12'h000;

			4858: dout = 12'h000;
			4859: dout = 12'h000;
			4860: dout = 12'h000;
			4861: dout = 12'h000;
			4862: dout = 12'h000;
			4863: dout = 12'h900;
			4864: dout = 12'hf10;
			4865: dout = 12'hf10;
			4866: dout = 12'hf10;
			4867: dout = 12'hf10;
			4868: dout = 12'hf10;
			4869: dout = 12'hf10;
			4870: dout = 12'hf10;
			4871: dout = 12'hf10;
			4872: dout = 12'hf10;
			4873: dout = 12'hf10;
			4874: dout = 12'hf10;
			4875: dout = 12'hf10;
			4876: dout = 12'hf10;
			4877: dout = 12'h100;
			4878: dout = 12'h000;
			4879: dout = 12'h000;
			4880: dout = 12'h000;
			4881: dout = 12'h600;
			4882: dout = 12'hf10;
			4883: dout = 12'hf10;
			4884: dout = 12'hf10;
			4885: dout = 12'hf10;
			4886: dout = 12'hf10;
			4887: dout = 12'hf10;
			4888: dout = 12'hf10;
			4889: dout = 12'h300;
			4890: dout = 12'h000;
			4891: dout = 12'h000;
			4892: dout = 12'h000;
			4893: dout = 12'h400;
			4894: dout = 12'hf10;
			4895: dout = 12'hf10;
			4896: dout = 12'hc10;
			4897: dout = 12'h000;
			4898: dout = 12'h000;
			4899: dout = 12'h000;
			4900: dout = 12'h000;
			4901: dout = 12'h000;
			4902: dout = 12'h000;
			4903: dout = 12'h000;
			4904: dout = 12'h000;
			4905: dout = 12'h200;
			4906: dout = 12'hf10;
			4907: dout = 12'hf10;
			4908: dout = 12'he10;
			4909: dout = 12'h000;
			4910: dout = 12'hb10;
			4911: dout = 12'hf10;
			4912: dout = 12'hf10;
			4913: dout = 12'hf10;
			4914: dout = 12'hf10;
			4915: dout = 12'hf10;
			4916: dout = 12'hf10;
			4917: dout = 12'hf10;
			4918: dout = 12'hf10;
			4919: dout = 12'hf10;
			4920: dout = 12'hf10;
			4921: dout = 12'hf10;
			4922: dout = 12'hf10;
			4923: dout = 12'hf10;
			4924: dout = 12'hf10;
			4925: dout = 12'h800;
			4926: dout = 12'h000;
			4927: dout = 12'h000;
			4928: dout = 12'h000;
			4929: dout = 12'h000;
			4930: dout = 12'h000;
			4931: dout = 12'h000;
			4932: dout = 12'h000;
			4933: dout = 12'h000;
			4934: dout = 12'h000;
			4935: dout = 12'h000;
			4936: dout = 12'h000;
			4937: dout = 12'h600;
			4938: dout = 12'hf10;
			4939: dout = 12'hf10;
			4940: dout = 12'hf10;
			4941: dout = 12'hf10;
			4942: dout = 12'hf10;
			4943: dout = 12'hf10;
			4944: dout = 12'hf10;
			4945: dout = 12'hf10;
			4946: dout = 12'hf10;
			4947: dout = 12'hf10;
			4948: dout = 12'hf10;
			4949: dout = 12'hc10;
			4950: dout = 12'h000;
			4951: dout = 12'h000;
			4952: dout = 12'h000;
			4953: dout = 12'h000;
			4954: dout = 12'he10;
			4955: dout = 12'hf10;
			4956: dout = 12'hf10;
			4957: dout = 12'h200;
			4958: dout = 12'h000;
			4959: dout = 12'h000;
			4960: dout = 12'h000;
			4961: dout = 12'h000;
			4962: dout = 12'h000;
			4963: dout = 12'h000;
			4964: dout = 12'h000;
			4965: dout = 12'h000;
			4966: dout = 12'hc10;
			4967: dout = 12'hf10;
			4968: dout = 12'hf10;
			4969: dout = 12'h400;
			4970: dout = 12'h100;
			4971: dout = 12'hf10;
			4972: dout = 12'hf10;
			4973: dout = 12'hf10;
			4974: dout = 12'hf10;
			4975: dout = 12'hf10;
			4976: dout = 12'hf10;
			4977: dout = 12'hf10;
			4978: dout = 12'hf10;
			4979: dout = 12'hf10;
			4980: dout = 12'hf10;
			4981: dout = 12'hf10;
			4982: dout = 12'hf10;
			4983: dout = 12'hf10;
			4984: dout = 12'hf10;
			4985: dout = 12'hf10;
			4986: dout = 12'h000;
			4987: dout = 12'h900;
			4988: dout = 12'hf10;
			4989: dout = 12'hf10;
			4990: dout = 12'hf10;
			4991: dout = 12'hf10;
			4992: dout = 12'hf10;
			4993: dout = 12'hf10;
			4994: dout = 12'hf10;
			4995: dout = 12'hf10;
			4996: dout = 12'hf10;
			4997: dout = 12'hf10;
			4998: dout = 12'hf10;
			4999: dout = 12'hf10;
			5000: dout = 12'hf10;
			5001: dout = 12'h100;
			5002: dout = 12'h000;
			5003: dout = 12'h000;
			5004: dout = 12'h000;
			5005: dout = 12'h000;
			5006: dout = 12'h000;
			5007: dout = 12'h000;

			5008: dout = 12'h000;
			5009: dout = 12'h000;
			5010: dout = 12'h000;
			5011: dout = 12'h000;
			5012: dout = 12'h000;
			5013: dout = 12'h810;
			5014: dout = 12'hf20;
			5015: dout = 12'hf20;
			5016: dout = 12'hf20;
			5017: dout = 12'hf20;
			5018: dout = 12'hf20;
			5019: dout = 12'hf20;
			5020: dout = 12'hf20;
			5021: dout = 12'hf20;
			5022: dout = 12'hf20;
			5023: dout = 12'hf20;
			5024: dout = 12'hf20;
			5025: dout = 12'hf20;
			5026: dout = 12'hf20;
			5027: dout = 12'h200;
			5028: dout = 12'h000;
			5029: dout = 12'h000;
			5030: dout = 12'h000;
			5031: dout = 12'h500;
			5032: dout = 12'hf20;
			5033: dout = 12'hf20;
			5034: dout = 12'hf20;
			5035: dout = 12'hf20;
			5036: dout = 12'hf20;
			5037: dout = 12'hf20;
			5038: dout = 12'hf20;
			5039: dout = 12'h200;
			5040: dout = 12'h000;
			5041: dout = 12'h000;
			5042: dout = 12'h000;
			5043: dout = 12'h400;
			5044: dout = 12'hf20;
			5045: dout = 12'hf20;
			5046: dout = 12'hc10;
			5047: dout = 12'h000;
			5048: dout = 12'h000;
			5049: dout = 12'h000;
			5050: dout = 12'h000;
			5051: dout = 12'h000;
			5052: dout = 12'h000;
			5053: dout = 12'h000;
			5054: dout = 12'h000;
			5055: dout = 12'h200;
			5056: dout = 12'hf20;
			5057: dout = 12'hf20;
			5058: dout = 12'he10;
			5059: dout = 12'h000;
			5060: dout = 12'ha10;
			5061: dout = 12'hf20;
			5062: dout = 12'hf20;
			5063: dout = 12'hf20;
			5064: dout = 12'hf20;
			5065: dout = 12'hf20;
			5066: dout = 12'hf20;
			5067: dout = 12'hf20;
			5068: dout = 12'hf20;
			5069: dout = 12'hf20;
			5070: dout = 12'hf20;
			5071: dout = 12'hf20;
			5072: dout = 12'hf20;
			5073: dout = 12'hf20;
			5074: dout = 12'hf20;
			5075: dout = 12'h810;
			5076: dout = 12'h000;
			5077: dout = 12'h000;
			5078: dout = 12'h000;
			5079: dout = 12'h000;
			5080: dout = 12'h000;
			5081: dout = 12'h000;
			5082: dout = 12'h000;
			5083: dout = 12'h000;
			5084: dout = 12'h000;
			5085: dout = 12'h000;
			5086: dout = 12'h000;
			5087: dout = 12'h600;
			5088: dout = 12'hf20;
			5089: dout = 12'hf20;
			5090: dout = 12'hf20;
			5091: dout = 12'hf20;
			5092: dout = 12'hf20;
			5093: dout = 12'hf20;
			5094: dout = 12'hf20;
			5095: dout = 12'hf20;
			5096: dout = 12'hf20;
			5097: dout = 12'hf20;
			5098: dout = 12'hf20;
			5099: dout = 12'hc10;
			5100: dout = 12'h000;
			5101: dout = 12'h000;
			5102: dout = 12'h000;
			5103: dout = 12'h000;
			5104: dout = 12'hd10;
			5105: dout = 12'hf20;
			5106: dout = 12'hf20;
			5107: dout = 12'h200;
			5108: dout = 12'h000;
			5109: dout = 12'h000;
			5110: dout = 12'h000;
			5111: dout = 12'h000;
			5112: dout = 12'h000;
			5113: dout = 12'h000;
			5114: dout = 12'h000;
			5115: dout = 12'h000;
			5116: dout = 12'hc10;
			5117: dout = 12'hf20;
			5118: dout = 12'hf20;
			5119: dout = 12'h400;
			5120: dout = 12'h100;
			5121: dout = 12'hf20;
			5122: dout = 12'hf20;
			5123: dout = 12'hf20;
			5124: dout = 12'hf20;
			5125: dout = 12'hf20;
			5126: dout = 12'hf20;
			5127: dout = 12'hf20;
			5128: dout = 12'hf20;
			5129: dout = 12'hf20;
			5130: dout = 12'hf20;
			5131: dout = 12'hf20;
			5132: dout = 12'hf20;
			5133: dout = 12'hf20;
			5134: dout = 12'hf20;
			5135: dout = 12'hf20;
			5136: dout = 12'h000;
			5137: dout = 12'h810;
			5138: dout = 12'hf20;
			5139: dout = 12'hf20;
			5140: dout = 12'hf20;
			5141: dout = 12'hf20;
			5142: dout = 12'hf20;
			5143: dout = 12'hf20;
			5144: dout = 12'hf20;
			5145: dout = 12'hf20;
			5146: dout = 12'hf20;
			5147: dout = 12'hf20;
			5148: dout = 12'hf20;
			5149: dout = 12'hf20;
			5150: dout = 12'hf20;
			5151: dout = 12'h100;
			5152: dout = 12'h000;
			5153: dout = 12'h000;
			5154: dout = 12'h000;
			5155: dout = 12'h000;
			5156: dout = 12'h000;
			5157: dout = 12'h000;

			5158: dout = 12'h000;
			5159: dout = 12'h000;
			5160: dout = 12'h910;
			5161: dout = 12'hd20;
			5162: dout = 12'hd20;
			5163: dout = 12'h700;
			5164: dout = 12'h100;
			5165: dout = 12'h200;
			5166: dout = 12'h200;
			5167: dout = 12'h200;
			5168: dout = 12'h200;
			5169: dout = 12'h200;
			5170: dout = 12'h200;
			5171: dout = 12'h200;
			5172: dout = 12'h200;
			5173: dout = 12'h200;
			5174: dout = 12'h200;
			5175: dout = 12'h200;
			5176: dout = 12'h200;
			5177: dout = 12'h000;
			5178: dout = 12'h600;
			5179: dout = 12'he20;
			5180: dout = 12'hd20;
			5181: dout = 12'h910;
			5182: dout = 12'h100;
			5183: dout = 12'h200;
			5184: dout = 12'h200;
			5185: dout = 12'h200;
			5186: dout = 12'h200;
			5187: dout = 12'h200;
			5188: dout = 12'h200;
			5189: dout = 12'hb10;
			5190: dout = 12'hd20;
			5191: dout = 12'he20;
			5192: dout = 12'h300;
			5193: dout = 12'h300;
			5194: dout = 12'hf30;
			5195: dout = 12'hf30;
			5196: dout = 12'he20;
			5197: dout = 12'hd20;
			5198: dout = 12'he20;
			5199: dout = 12'hc10;
			5200: dout = 12'h000;
			5201: dout = 12'h000;
			5202: dout = 12'h300;
			5203: dout = 12'he20;
			5204: dout = 12'hd20;
			5205: dout = 12'hd20;
			5206: dout = 12'hf30;
			5207: dout = 12'hf30;
			5208: dout = 12'he20;
			5209: dout = 12'h000;
			5210: dout = 12'ha10;
			5211: dout = 12'hf30;
			5212: dout = 12'hf30;
			5213: dout = 12'h600;
			5214: dout = 12'h100;
			5215: dout = 12'h200;
			5216: dout = 12'h200;
			5217: dout = 12'h200;
			5218: dout = 12'h200;
			5219: dout = 12'h200;
			5220: dout = 12'h200;
			5221: dout = 12'h200;
			5222: dout = 12'h200;
			5223: dout = 12'h200;
			5224: dout = 12'h200;
			5225: dout = 12'h200;
			5226: dout = 12'h000;
			5227: dout = 12'h000;
			5228: dout = 12'h000;
			5229: dout = 12'h000;
			5230: dout = 12'h000;
			5231: dout = 12'h000;
			5232: dout = 12'h000;
			5233: dout = 12'h000;
			5234: dout = 12'h600;
			5235: dout = 12'he20;
			5236: dout = 12'hd20;
			5237: dout = 12'h910;
			5238: dout = 12'h100;
			5239: dout = 12'h200;
			5240: dout = 12'h200;
			5241: dout = 12'h200;
			5242: dout = 12'h200;
			5243: dout = 12'h200;
			5244: dout = 12'h200;
			5245: dout = 12'h200;
			5246: dout = 12'h200;
			5247: dout = 12'h200;
			5248: dout = 12'h200;
			5249: dout = 12'h500;
			5250: dout = 12'he20;
			5251: dout = 12'hd20;
			5252: dout = 12'hb10;
			5253: dout = 12'h000;
			5254: dout = 12'hd20;
			5255: dout = 12'hf30;
			5256: dout = 12'hf30;
			5257: dout = 12'h200;
			5258: dout = 12'h000;
			5259: dout = 12'h000;
			5260: dout = 12'h000;
			5261: dout = 12'h000;
			5262: dout = 12'h000;
			5263: dout = 12'h000;
			5264: dout = 12'h000;
			5265: dout = 12'h000;
			5266: dout = 12'hc20;
			5267: dout = 12'hf30;
			5268: dout = 12'hf30;
			5269: dout = 12'h400;
			5270: dout = 12'h100;
			5271: dout = 12'hf30;
			5272: dout = 12'hf30;
			5273: dout = 12'hd20;
			5274: dout = 12'h200;
			5275: dout = 12'h200;
			5276: dout = 12'h200;
			5277: dout = 12'h200;
			5278: dout = 12'h200;
			5279: dout = 12'h200;
			5280: dout = 12'h200;
			5281: dout = 12'h200;
			5282: dout = 12'h200;
			5283: dout = 12'h200;
			5284: dout = 12'h200;
			5285: dout = 12'h300;
			5286: dout = 12'h000;
			5287: dout = 12'h910;
			5288: dout = 12'hf30;
			5289: dout = 12'hf30;
			5290: dout = 12'h810;
			5291: dout = 12'h100;
			5292: dout = 12'h200;
			5293: dout = 12'h200;
			5294: dout = 12'h200;
			5295: dout = 12'h200;
			5296: dout = 12'h200;
			5297: dout = 12'h200;
			5298: dout = 12'h200;
			5299: dout = 12'h200;
			5300: dout = 12'h200;
			5301: dout = 12'hc20;
			5302: dout = 12'he20;
			5303: dout = 12'he20;
			5304: dout = 12'h200;
			5305: dout = 12'h000;
			5306: dout = 12'h000;
			5307: dout = 12'h000;

			5308: dout = 12'h000;
			5309: dout = 12'h000;
			5310: dout = 12'h910;
			5311: dout = 12'hf40;
			5312: dout = 12'hf40;
			5313: dout = 12'h710;
			5314: dout = 12'h000;
			5315: dout = 12'h000;
			5316: dout = 12'h000;
			5317: dout = 12'h000;
			5318: dout = 12'h000;
			5319: dout = 12'h000;
			5320: dout = 12'h000;
			5321: dout = 12'h000;
			5322: dout = 12'h000;
			5323: dout = 12'h000;
			5324: dout = 12'h000;
			5325: dout = 12'h000;
			5326: dout = 12'h000;
			5327: dout = 12'h000;
			5328: dout = 12'h600;
			5329: dout = 12'hf40;
			5330: dout = 12'hf40;
			5331: dout = 12'ha20;
			5332: dout = 12'h000;
			5333: dout = 12'h000;
			5334: dout = 12'h000;
			5335: dout = 12'h000;
			5336: dout = 12'h000;
			5337: dout = 12'h000;
			5338: dout = 12'h000;
			5339: dout = 12'hd20;
			5340: dout = 12'hf40;
			5341: dout = 12'hf40;
			5342: dout = 12'h200;
			5343: dout = 12'h300;
			5344: dout = 12'hf40;
			5345: dout = 12'hf40;
			5346: dout = 12'hf40;
			5347: dout = 12'hf40;
			5348: dout = 12'hf40;
			5349: dout = 12'hd20;
			5350: dout = 12'h000;
			5351: dout = 12'h000;
			5352: dout = 12'h300;
			5353: dout = 12'hf40;
			5354: dout = 12'hf40;
			5355: dout = 12'hf40;
			5356: dout = 12'hf40;
			5357: dout = 12'hf40;
			5358: dout = 12'he30;
			5359: dout = 12'h000;
			5360: dout = 12'ha20;
			5361: dout = 12'hf40;
			5362: dout = 12'hf40;
			5363: dout = 12'h500;
			5364: dout = 12'h000;
			5365: dout = 12'h000;
			5366: dout = 12'h000;
			5367: dout = 12'h000;
			5368: dout = 12'h000;
			5369: dout = 12'h000;
			5370: dout = 12'h000;
			5371: dout = 12'h000;
			5372: dout = 12'h000;
			5373: dout = 12'h000;
			5374: dout = 12'h000;
			5375: dout = 12'h000;
			5376: dout = 12'h000;
			5377: dout = 12'h000;
			5378: dout = 12'h000;
			5379: dout = 12'h000;
			5380: dout = 12'h000;
			5381: dout = 12'h000;
			5382: dout = 12'h000;
			5383: dout = 12'h000;
			5384: dout = 12'h710;
			5385: dout = 12'hf40;
			5386: dout = 12'hf40;
			5387: dout = 12'h910;
			5388: dout = 12'h000;
			5389: dout = 12'h000;
			5390: dout = 12'h000;
			5391: dout = 12'h000;
			5392: dout = 12'h000;
			5393: dout = 12'h000;
			5394: dout = 12'h000;
			5395: dout = 12'h000;
			5396: dout = 12'h000;
			5397: dout = 12'h000;
			5398: dout = 12'h000;
			5399: dout = 12'h400;
			5400: dout = 12'hf40;
			5401: dout = 12'hf40;
			5402: dout = 12'hc20;
			5403: dout = 12'h000;
			5404: dout = 12'hd30;
			5405: dout = 12'hf40;
			5406: dout = 12'hf40;
			5407: dout = 12'h200;
			5408: dout = 12'h000;
			5409: dout = 12'h000;
			5410: dout = 12'h000;
			5411: dout = 12'h000;
			5412: dout = 12'h000;
			5413: dout = 12'h000;
			5414: dout = 12'h000;
			5415: dout = 12'h000;
			5416: dout = 12'hc20;
			5417: dout = 12'hf40;
			5418: dout = 12'hf40;
			5419: dout = 12'h400;
			5420: dout = 12'h100;
			5421: dout = 12'hf40;
			5422: dout = 12'hf40;
			5423: dout = 12'he30;
			5424: dout = 12'h000;
			5425: dout = 12'h000;
			5426: dout = 12'h000;
			5427: dout = 12'h000;
			5428: dout = 12'h000;
			5429: dout = 12'h000;
			5430: dout = 12'h000;
			5431: dout = 12'h000;
			5432: dout = 12'h000;
			5433: dout = 12'h000;
			5434: dout = 12'h000;
			5435: dout = 12'h000;
			5436: dout = 12'h000;
			5437: dout = 12'h910;
			5438: dout = 12'hf40;
			5439: dout = 12'hf40;
			5440: dout = 12'h710;
			5441: dout = 12'h000;
			5442: dout = 12'h000;
			5443: dout = 12'h000;
			5444: dout = 12'h000;
			5445: dout = 12'h000;
			5446: dout = 12'h000;
			5447: dout = 12'h000;
			5448: dout = 12'h000;
			5449: dout = 12'h000;
			5450: dout = 12'h000;
			5451: dout = 12'he30;
			5452: dout = 12'hf40;
			5453: dout = 12'hf40;
			5454: dout = 12'h200;
			5455: dout = 12'h000;
			5456: dout = 12'h000;
			5457: dout = 12'h000;

			5458: dout = 12'h000;
			5459: dout = 12'h000;
			5460: dout = 12'h920;
			5461: dout = 12'hf50;
			5462: dout = 12'hf50;
			5463: dout = 12'h710;
			5464: dout = 12'h000;
			5465: dout = 12'h000;
			5466: dout = 12'h000;
			5467: dout = 12'h000;
			5468: dout = 12'h000;
			5469: dout = 12'h000;
			5470: dout = 12'h000;
			5471: dout = 12'h000;
			5472: dout = 12'h000;
			5473: dout = 12'h000;
			5474: dout = 12'h000;
			5475: dout = 12'h000;
			5476: dout = 12'h000;
			5477: dout = 12'h000;
			5478: dout = 12'h610;
			5479: dout = 12'hf50;
			5480: dout = 12'hf50;
			5481: dout = 12'ha20;
			5482: dout = 12'h000;
			5483: dout = 12'h000;
			5484: dout = 12'h000;
			5485: dout = 12'h000;
			5486: dout = 12'h000;
			5487: dout = 12'h000;
			5488: dout = 12'h000;
			5489: dout = 12'hd30;
			5490: dout = 12'hf50;
			5491: dout = 12'hf50;
			5492: dout = 12'h200;
			5493: dout = 12'h300;
			5494: dout = 12'hf50;
			5495: dout = 12'hf50;
			5496: dout = 12'hf50;
			5497: dout = 12'hf40;
			5498: dout = 12'hf50;
			5499: dout = 12'hc30;
			5500: dout = 12'h000;
			5501: dout = 12'h000;
			5502: dout = 12'h200;
			5503: dout = 12'hf50;
			5504: dout = 12'hf50;
			5505: dout = 12'hf40;
			5506: dout = 12'hf50;
			5507: dout = 12'hf50;
			5508: dout = 12'he30;
			5509: dout = 12'h000;
			5510: dout = 12'ha20;
			5511: dout = 12'hf50;
			5512: dout = 12'hf50;
			5513: dout = 12'h500;
			5514: dout = 12'h000;
			5515: dout = 12'h000;
			5516: dout = 12'h000;
			5517: dout = 12'h000;
			5518: dout = 12'h000;
			5519: dout = 12'h000;
			5520: dout = 12'h000;
			5521: dout = 12'h000;
			5522: dout = 12'h000;
			5523: dout = 12'h000;
			5524: dout = 12'h000;
			5525: dout = 12'h000;
			5526: dout = 12'h000;
			5527: dout = 12'h000;
			5528: dout = 12'h000;
			5529: dout = 12'h000;
			5530: dout = 12'h000;
			5531: dout = 12'h000;
			5532: dout = 12'h000;
			5533: dout = 12'h000;
			5534: dout = 12'h710;
			5535: dout = 12'hf50;
			5536: dout = 12'hf50;
			5537: dout = 12'h920;
			5538: dout = 12'h000;
			5539: dout = 12'h000;
			5540: dout = 12'h000;
			5541: dout = 12'h000;
			5542: dout = 12'h000;
			5543: dout = 12'h000;
			5544: dout = 12'h000;
			5545: dout = 12'h000;
			5546: dout = 12'h000;
			5547: dout = 12'h000;
			5548: dout = 12'h000;
			5549: dout = 12'h400;
			5550: dout = 12'hf50;
			5551: dout = 12'hf50;
			5552: dout = 12'hc20;
			5553: dout = 12'h000;
			5554: dout = 12'hd30;
			5555: dout = 12'hf50;
			5556: dout = 12'hf50;
			5557: dout = 12'h200;
			5558: dout = 12'h000;
			5559: dout = 12'h000;
			5560: dout = 12'h000;
			5561: dout = 12'h000;
			5562: dout = 12'h000;
			5563: dout = 12'h000;
			5564: dout = 12'h000;
			5565: dout = 12'h000;
			5566: dout = 12'hc20;
			5567: dout = 12'hf50;
			5568: dout = 12'hf50;
			5569: dout = 12'h400;
			5570: dout = 12'h100;
			5571: dout = 12'hf50;
			5572: dout = 12'hf50;
			5573: dout = 12'hd30;
			5574: dout = 12'h000;
			5575: dout = 12'h000;
			5576: dout = 12'h000;
			5577: dout = 12'h000;
			5578: dout = 12'h000;
			5579: dout = 12'h000;
			5580: dout = 12'h000;
			5581: dout = 12'h000;
			5582: dout = 12'h000;
			5583: dout = 12'h000;
			5584: dout = 12'h000;
			5585: dout = 12'h000;
			5586: dout = 12'h000;
			5587: dout = 12'h910;
			5588: dout = 12'hf50;
			5589: dout = 12'hf50;
			5590: dout = 12'h710;
			5591: dout = 12'h000;
			5592: dout = 12'h000;
			5593: dout = 12'h000;
			5594: dout = 12'h000;
			5595: dout = 12'h000;
			5596: dout = 12'h000;
			5597: dout = 12'h000;
			5598: dout = 12'h000;
			5599: dout = 12'h000;
			5600: dout = 12'h000;
			5601: dout = 12'he30;
			5602: dout = 12'hf50;
			5603: dout = 12'hf40;
			5604: dout = 12'h200;
			5605: dout = 12'h000;
			5606: dout = 12'h000;
			5607: dout = 12'h000;

			5608: dout = 12'h000;
			5609: dout = 12'h000;
			5610: dout = 12'h920;
			5611: dout = 12'hf60;
			5612: dout = 12'hf60;
			5613: dout = 12'h710;
			5614: dout = 12'h000;
			5615: dout = 12'h000;
			5616: dout = 12'h000;
			5617: dout = 12'h000;
			5618: dout = 12'h000;
			5619: dout = 12'h000;
			5620: dout = 12'h000;
			5621: dout = 12'hd30;
			5622: dout = 12'hd40;
			5623: dout = 12'hd30;
			5624: dout = 12'hd30;
			5625: dout = 12'hd40;
			5626: dout = 12'hd30;
			5627: dout = 12'h100;
			5628: dout = 12'h610;
			5629: dout = 12'hf60;
			5630: dout = 12'hf60;
			5631: dout = 12'hd40;
			5632: dout = 12'hd30;
			5633: dout = 12'hd30;
			5634: dout = 12'hd30;
			5635: dout = 12'hd30;
			5636: dout = 12'hd30;
			5637: dout = 12'hd30;
			5638: dout = 12'hc30;
			5639: dout = 12'he50;
			5640: dout = 12'hf60;
			5641: dout = 12'hf60;
			5642: dout = 12'h200;
			5643: dout = 12'h300;
			5644: dout = 12'hf60;
			5645: dout = 12'hf60;
			5646: dout = 12'hb30;
			5647: dout = 12'h000;
			5648: dout = 12'h000;
			5649: dout = 12'h400;
			5650: dout = 12'hd40;
			5651: dout = 12'hd40;
			5652: dout = 12'hb20;
			5653: dout = 12'h000;
			5654: dout = 12'h000;
			5655: dout = 12'h300;
			5656: dout = 12'hf60;
			5657: dout = 12'hf60;
			5658: dout = 12'he40;
			5659: dout = 12'h000;
			5660: dout = 12'ha20;
			5661: dout = 12'hf60;
			5662: dout = 12'hf60;
			5663: dout = 12'hd40;
			5664: dout = 12'hd30;
			5665: dout = 12'hd30;
			5666: dout = 12'hd40;
			5667: dout = 12'hc30;
			5668: dout = 12'h000;
			5669: dout = 12'h000;
			5670: dout = 12'h000;
			5671: dout = 12'h000;
			5672: dout = 12'h000;
			5673: dout = 12'h000;
			5674: dout = 12'h000;
			5675: dout = 12'h000;
			5676: dout = 12'h000;
			5677: dout = 12'h000;
			5678: dout = 12'h000;
			5679: dout = 12'h000;
			5680: dout = 12'h000;
			5681: dout = 12'h000;
			5682: dout = 12'h000;
			5683: dout = 12'h000;
			5684: dout = 12'h710;
			5685: dout = 12'hf60;
			5686: dout = 12'hf60;
			5687: dout = 12'h920;
			5688: dout = 12'h000;
			5689: dout = 12'h000;
			5690: dout = 12'h000;
			5691: dout = 12'h000;
			5692: dout = 12'h000;
			5693: dout = 12'h000;
			5694: dout = 12'h000;
			5695: dout = 12'h000;
			5696: dout = 12'h000;
			5697: dout = 12'h000;
			5698: dout = 12'h000;
			5699: dout = 12'h400;
			5700: dout = 12'hf60;
			5701: dout = 12'hf60;
			5702: dout = 12'hc30;
			5703: dout = 12'h000;
			5704: dout = 12'he40;
			5705: dout = 12'hf70;
			5706: dout = 12'hf70;
			5707: dout = 12'h200;
			5708: dout = 12'h000;
			5709: dout = 12'h000;
			5710: dout = 12'h000;
			5711: dout = 12'h000;
			5712: dout = 12'h000;
			5713: dout = 12'h000;
			5714: dout = 12'h000;
			5715: dout = 12'h000;
			5716: dout = 12'hc30;
			5717: dout = 12'hf70;
			5718: dout = 12'hf70;
			5719: dout = 12'h400;
			5720: dout = 12'h100;
			5721: dout = 12'hf60;
			5722: dout = 12'hf60;
			5723: dout = 12'he50;
			5724: dout = 12'hc30;
			5725: dout = 12'hd30;
			5726: dout = 12'hd30;
			5727: dout = 12'he40;
			5728: dout = 12'h600;
			5729: dout = 12'h000;
			5730: dout = 12'h000;
			5731: dout = 12'h000;
			5732: dout = 12'h000;
			5733: dout = 12'h000;
			5734: dout = 12'h000;
			5735: dout = 12'h000;
			5736: dout = 12'h000;
			5737: dout = 12'h920;
			5738: dout = 12'hf60;
			5739: dout = 12'hf60;
			5740: dout = 12'hd40;
			5741: dout = 12'hd30;
			5742: dout = 12'hd30;
			5743: dout = 12'hd30;
			5744: dout = 12'hd30;
			5745: dout = 12'hd30;
			5746: dout = 12'hd30;
			5747: dout = 12'hd30;
			5748: dout = 12'hd30;
			5749: dout = 12'hd40;
			5750: dout = 12'hd30;
			5751: dout = 12'h300;
			5752: dout = 12'h100;
			5753: dout = 12'h100;
			5754: dout = 12'h000;
			5755: dout = 12'h000;
			5756: dout = 12'h000;
			5757: dout = 12'h000;

			5758: dout = 12'h000;
			5759: dout = 12'h000;
			5760: dout = 12'h920;
			5761: dout = 12'hf70;
			5762: dout = 12'hf70;
			5763: dout = 12'h710;
			5764: dout = 12'h000;
			5765: dout = 12'h000;
			5766: dout = 12'h000;
			5767: dout = 12'h000;
			5768: dout = 12'h000;
			5769: dout = 12'h000;
			5770: dout = 12'h000;
			5771: dout = 12'hf50;
			5772: dout = 12'hf70;
			5773: dout = 12'hf70;
			5774: dout = 12'hf70;
			5775: dout = 12'hf70;
			5776: dout = 12'hf60;
			5777: dout = 12'h100;
			5778: dout = 12'h610;
			5779: dout = 12'hf70;
			5780: dout = 12'hf70;
			5781: dout = 12'hf70;
			5782: dout = 12'hf70;
			5783: dout = 12'hf70;
			5784: dout = 12'hf70;
			5785: dout = 12'hf70;
			5786: dout = 12'hf70;
			5787: dout = 12'hf70;
			5788: dout = 12'hf70;
			5789: dout = 12'hf70;
			5790: dout = 12'hf70;
			5791: dout = 12'hf70;
			5792: dout = 12'h200;
			5793: dout = 12'h300;
			5794: dout = 12'hf70;
			5795: dout = 12'hf70;
			5796: dout = 12'hc40;
			5797: dout = 12'h000;
			5798: dout = 12'h000;
			5799: dout = 12'h300;
			5800: dout = 12'hf70;
			5801: dout = 12'hf70;
			5802: dout = 12'hd40;
			5803: dout = 12'h000;
			5804: dout = 12'h000;
			5805: dout = 12'h200;
			5806: dout = 12'hf70;
			5807: dout = 12'hf70;
			5808: dout = 12'he40;
			5809: dout = 12'h000;
			5810: dout = 12'ha30;
			5811: dout = 12'hf70;
			5812: dout = 12'hf70;
			5813: dout = 12'hf70;
			5814: dout = 12'hf70;
			5815: dout = 12'hf70;
			5816: dout = 12'hf70;
			5817: dout = 12'hf50;
			5818: dout = 12'h000;
			5819: dout = 12'h000;
			5820: dout = 12'h000;
			5821: dout = 12'h000;
			5822: dout = 12'h000;
			5823: dout = 12'h000;
			5824: dout = 12'h000;
			5825: dout = 12'h000;
			5826: dout = 12'h000;
			5827: dout = 12'h000;
			5828: dout = 12'h000;
			5829: dout = 12'h000;
			5830: dout = 12'h000;
			5831: dout = 12'h000;
			5832: dout = 12'h000;
			5833: dout = 12'h000;
			5834: dout = 12'h710;
			5835: dout = 12'hf70;
			5836: dout = 12'hf70;
			5837: dout = 12'h920;
			5838: dout = 12'h000;
			5839: dout = 12'h000;
			5840: dout = 12'h000;
			5841: dout = 12'h000;
			5842: dout = 12'h000;
			5843: dout = 12'h000;
			5844: dout = 12'h000;
			5845: dout = 12'h000;
			5846: dout = 12'h000;
			5847: dout = 12'h000;
			5848: dout = 12'h000;
			5849: dout = 12'h400;
			5850: dout = 12'hf70;
			5851: dout = 12'hf70;
			5852: dout = 12'hc30;
			5853: dout = 12'h000;
			5854: dout = 12'h810;
			5855: dout = 12'h820;
			5856: dout = 12'h820;
			5857: dout = 12'h700;
			5858: dout = 12'h610;
			5859: dout = 12'h610;
			5860: dout = 12'h200;
			5861: dout = 12'h000;
			5862: dout = 12'h000;
			5863: dout = 12'h600;
			5864: dout = 12'h610;
			5865: dout = 12'h610;
			5866: dout = 12'h810;
			5867: dout = 12'h820;
			5868: dout = 12'h920;
			5869: dout = 12'h300;
			5870: dout = 12'h200;
			5871: dout = 12'hf70;
			5872: dout = 12'hf70;
			5873: dout = 12'hf70;
			5874: dout = 12'hf70;
			5875: dout = 12'hf70;
			5876: dout = 12'hf70;
			5877: dout = 12'hf80;
			5878: dout = 12'h610;
			5879: dout = 12'h000;
			5880: dout = 12'h000;
			5881: dout = 12'h000;
			5882: dout = 12'h000;
			5883: dout = 12'h000;
			5884: dout = 12'h000;
			5885: dout = 12'h000;
			5886: dout = 12'h000;
			5887: dout = 12'h920;
			5888: dout = 12'hf70;
			5889: dout = 12'hf70;
			5890: dout = 12'hf70;
			5891: dout = 12'hf70;
			5892: dout = 12'hf70;
			5893: dout = 12'hf70;
			5894: dout = 12'hf70;
			5895: dout = 12'hf70;
			5896: dout = 12'hf70;
			5897: dout = 12'hf70;
			5898: dout = 12'hf70;
			5899: dout = 12'hf70;
			5900: dout = 12'hf60;
			5901: dout = 12'h100;
			5902: dout = 12'h000;
			5903: dout = 12'h000;
			5904: dout = 12'h000;
			5905: dout = 12'h000;
			5906: dout = 12'h000;
			5907: dout = 12'h000;

			5908: dout = 12'h000;
			5909: dout = 12'h000;
			5910: dout = 12'h920;
			5911: dout = 12'hf80;
			5912: dout = 12'hf80;
			5913: dout = 12'h710;
			5914: dout = 12'h000;
			5915: dout = 12'h000;
			5916: dout = 12'h000;
			5917: dout = 12'h000;
			5918: dout = 12'h000;
			5919: dout = 12'h000;
			5920: dout = 12'h000;
			5921: dout = 12'hf60;
			5922: dout = 12'hf80;
			5923: dout = 12'hf70;
			5924: dout = 12'hf80;
			5925: dout = 12'hf80;
			5926: dout = 12'hf70;
			5927: dout = 12'h100;
			5928: dout = 12'h610;
			5929: dout = 12'hf80;
			5930: dout = 12'hf80;
			5931: dout = 12'hf80;
			5932: dout = 12'hf80;
			5933: dout = 12'hf80;
			5934: dout = 12'hf80;
			5935: dout = 12'hf80;
			5936: dout = 12'hf80;
			5937: dout = 12'hf80;
			5938: dout = 12'hf80;
			5939: dout = 12'hf80;
			5940: dout = 12'hf80;
			5941: dout = 12'hf80;
			5942: dout = 12'h200;
			5943: dout = 12'h300;
			5944: dout = 12'hf80;
			5945: dout = 12'hf80;
			5946: dout = 12'hc40;
			5947: dout = 12'h000;
			5948: dout = 12'h000;
			5949: dout = 12'h300;
			5950: dout = 12'hf80;
			5951: dout = 12'hf80;
			5952: dout = 12'hd50;
			5953: dout = 12'h000;
			5954: dout = 12'h000;
			5955: dout = 12'h200;
			5956: dout = 12'hf80;
			5957: dout = 12'hf80;
			5958: dout = 12'he50;
			5959: dout = 12'h000;
			5960: dout = 12'ha30;
			5961: dout = 12'hf80;
			5962: dout = 12'hf80;
			5963: dout = 12'hf80;
			5964: dout = 12'hf80;
			5965: dout = 12'hf80;
			5966: dout = 12'hf80;
			5967: dout = 12'hf60;
			5968: dout = 12'h000;
			5969: dout = 12'h000;
			5970: dout = 12'h000;
			5971: dout = 12'h000;
			5972: dout = 12'h000;
			5973: dout = 12'h000;
			5974: dout = 12'h000;
			5975: dout = 12'h000;
			5976: dout = 12'h000;
			5977: dout = 12'h000;
			5978: dout = 12'h000;
			5979: dout = 12'h000;
			5980: dout = 12'h000;
			5981: dout = 12'h000;
			5982: dout = 12'h000;
			5983: dout = 12'h000;
			5984: dout = 12'h710;
			5985: dout = 12'hf80;
			5986: dout = 12'hf80;
			5987: dout = 12'h920;
			5988: dout = 12'h000;
			5989: dout = 12'h000;
			5990: dout = 12'h000;
			5991: dout = 12'h000;
			5992: dout = 12'h000;
			5993: dout = 12'h000;
			5994: dout = 12'h000;
			5995: dout = 12'h000;
			5996: dout = 12'h000;
			5997: dout = 12'h000;
			5998: dout = 12'h000;
			5999: dout = 12'h400;
			6000: dout = 12'hf80;
			6001: dout = 12'hf80;
			6002: dout = 12'hc40;
			6003: dout = 12'h000;
			6004: dout = 12'h000;
			6005: dout = 12'h000;
			6006: dout = 12'h000;
			6007: dout = 12'he50;
			6008: dout = 12'hf90;
			6009: dout = 12'hf90;
			6010: dout = 12'h300;
			6011: dout = 12'h000;
			6012: dout = 12'h000;
			6013: dout = 12'hd40;
			6014: dout = 12'hf90;
			6015: dout = 12'hf90;
			6016: dout = 12'h300;
			6017: dout = 12'h000;
			6018: dout = 12'h000;
			6019: dout = 12'h000;
			6020: dout = 12'h200;
			6021: dout = 12'hf80;
			6022: dout = 12'hf80;
			6023: dout = 12'hf80;
			6024: dout = 12'hf80;
			6025: dout = 12'hf80;
			6026: dout = 12'hf80;
			6027: dout = 12'hf80;
			6028: dout = 12'h610;
			6029: dout = 12'h000;
			6030: dout = 12'h000;
			6031: dout = 12'h000;
			6032: dout = 12'h000;
			6033: dout = 12'h000;
			6034: dout = 12'h000;
			6035: dout = 12'h000;
			6036: dout = 12'h000;
			6037: dout = 12'h920;
			6038: dout = 12'hf80;
			6039: dout = 12'hf80;
			6040: dout = 12'hf80;
			6041: dout = 12'hf80;
			6042: dout = 12'hf80;
			6043: dout = 12'hf80;
			6044: dout = 12'hf80;
			6045: dout = 12'hf80;
			6046: dout = 12'hf80;
			6047: dout = 12'hf80;
			6048: dout = 12'hf80;
			6049: dout = 12'hf80;
			6050: dout = 12'hf70;
			6051: dout = 12'h200;
			6052: dout = 12'h000;
			6053: dout = 12'h000;
			6054: dout = 12'h000;
			6055: dout = 12'h000;
			6056: dout = 12'h000;
			6057: dout = 12'h000;

			6058: dout = 12'h000;
			6059: dout = 12'h000;
			6060: dout = 12'h930;
			6061: dout = 12'hf90;
			6062: dout = 12'hf90;
			6063: dout = 12'h720;
			6064: dout = 12'h000;
			6065: dout = 12'h000;
			6066: dout = 12'h000;
			6067: dout = 12'h000;
			6068: dout = 12'h000;
			6069: dout = 12'h000;
			6070: dout = 12'h000;
			6071: dout = 12'h200;
			6072: dout = 12'h200;
			6073: dout = 12'h200;
			6074: dout = 12'hd60;
			6075: dout = 12'hf90;
			6076: dout = 12'hf80;
			6077: dout = 12'h100;
			6078: dout = 12'h610;
			6079: dout = 12'hf90;
			6080: dout = 12'hf90;
			6081: dout = 12'ha30;
			6082: dout = 12'h100;
			6083: dout = 12'h200;
			6084: dout = 12'h200;
			6085: dout = 12'h200;
			6086: dout = 12'h200;
			6087: dout = 12'h200;
			6088: dout = 12'h100;
			6089: dout = 12'hc50;
			6090: dout = 12'hf90;
			6091: dout = 12'hf90;
			6092: dout = 12'h200;
			6093: dout = 12'h300;
			6094: dout = 12'hf90;
			6095: dout = 12'hf90;
			6096: dout = 12'hc40;
			6097: dout = 12'h000;
			6098: dout = 12'h000;
			6099: dout = 12'h100;
			6100: dout = 12'h200;
			6101: dout = 12'h200;
			6102: dout = 12'h200;
			6103: dout = 12'h000;
			6104: dout = 12'h000;
			6105: dout = 12'h200;
			6106: dout = 12'hf90;
			6107: dout = 12'hf90;
			6108: dout = 12'he50;
			6109: dout = 12'h000;
			6110: dout = 12'ha30;
			6111: dout = 12'hf90;
			6112: dout = 12'hf90;
			6113: dout = 12'h600;
			6114: dout = 12'h100;
			6115: dout = 12'h200;
			6116: dout = 12'h200;
			6117: dout = 12'h200;
			6118: dout = 12'h000;
			6119: dout = 12'h000;
			6120: dout = 12'h000;
			6121: dout = 12'h000;
			6122: dout = 12'h000;
			6123: dout = 12'h000;
			6124: dout = 12'h000;
			6125: dout = 12'h000;
			6126: dout = 12'h000;
			6127: dout = 12'h000;
			6128: dout = 12'h000;
			6129: dout = 12'h000;
			6130: dout = 12'h000;
			6131: dout = 12'h000;
			6132: dout = 12'h000;
			6133: dout = 12'h000;
			6134: dout = 12'h710;
			6135: dout = 12'hf90;
			6136: dout = 12'hf90;
			6137: dout = 12'h930;
			6138: dout = 12'h000;
			6139: dout = 12'h000;
			6140: dout = 12'h000;
			6141: dout = 12'h000;
			6142: dout = 12'h000;
			6143: dout = 12'h000;
			6144: dout = 12'h000;
			6145: dout = 12'h000;
			6146: dout = 12'h000;
			6147: dout = 12'h000;
			6148: dout = 12'h000;
			6149: dout = 12'h400;
			6150: dout = 12'hf90;
			6151: dout = 12'hf90;
			6152: dout = 12'hc40;
			6153: dout = 12'h000;
			6154: dout = 12'h000;
			6155: dout = 12'h000;
			6156: dout = 12'h000;
			6157: dout = 12'hd50;
			6158: dout = 12'hf90;
			6159: dout = 12'hf90;
			6160: dout = 12'h300;
			6161: dout = 12'h000;
			6162: dout = 12'h000;
			6163: dout = 12'hc50;
			6164: dout = 12'hf90;
			6165: dout = 12'hf90;
			6166: dout = 12'h400;
			6167: dout = 12'h000;
			6168: dout = 12'h000;
			6169: dout = 12'h000;
			6170: dout = 12'h200;
			6171: dout = 12'hf80;
			6172: dout = 12'hf90;
			6173: dout = 12'hd50;
			6174: dout = 12'h100;
			6175: dout = 12'h200;
			6176: dout = 12'h200;
			6177: dout = 12'h200;
			6178: dout = 12'h100;
			6179: dout = 12'h000;
			6180: dout = 12'h000;
			6181: dout = 12'h000;
			6182: dout = 12'h000;
			6183: dout = 12'h000;
			6184: dout = 12'h000;
			6185: dout = 12'h000;
			6186: dout = 12'h000;
			6187: dout = 12'h920;
			6188: dout = 12'hf90;
			6189: dout = 12'hf90;
			6190: dout = 12'h710;
			6191: dout = 12'h100;
			6192: dout = 12'h200;
			6193: dout = 12'h200;
			6194: dout = 12'h200;
			6195: dout = 12'h100;
			6196: dout = 12'h710;
			6197: dout = 12'hf90;
			6198: dout = 12'hf90;
			6199: dout = 12'h920;
			6200: dout = 12'h100;
			6201: dout = 12'h000;
			6202: dout = 12'h000;
			6203: dout = 12'h000;
			6204: dout = 12'h000;
			6205: dout = 12'h000;
			6206: dout = 12'h000;
			6207: dout = 12'h000;

			6208: dout = 12'h000;
			6209: dout = 12'h000;
			6210: dout = 12'h930;
			6211: dout = 12'hfa0;
			6212: dout = 12'hfa0;
			6213: dout = 12'h720;
			6214: dout = 12'h000;
			6215: dout = 12'h000;
			6216: dout = 12'h000;
			6217: dout = 12'h000;
			6218: dout = 12'h000;
			6219: dout = 12'h000;
			6220: dout = 12'h000;
			6221: dout = 12'h000;
			6222: dout = 12'h000;
			6223: dout = 12'h000;
			6224: dout = 12'he70;
			6225: dout = 12'hfa0;
			6226: dout = 12'hf90;
			6227: dout = 12'h100;
			6228: dout = 12'h610;
			6229: dout = 12'hfa0;
			6230: dout = 12'hfa0;
			6231: dout = 12'ha30;
			6232: dout = 12'h000;
			6233: dout = 12'h000;
			6234: dout = 12'h000;
			6235: dout = 12'h000;
			6236: dout = 12'h000;
			6237: dout = 12'h000;
			6238: dout = 12'h000;
			6239: dout = 12'hd60;
			6240: dout = 12'hfa0;
			6241: dout = 12'hfa0;
			6242: dout = 12'h200;
			6243: dout = 12'h300;
			6244: dout = 12'hfa0;
			6245: dout = 12'hfa0;
			6246: dout = 12'hc50;
			6247: dout = 12'h000;
			6248: dout = 12'h000;
			6249: dout = 12'h000;
			6250: dout = 12'h000;
			6251: dout = 12'h000;
			6252: dout = 12'h000;
			6253: dout = 12'h000;
			6254: dout = 12'h000;
			6255: dout = 12'h200;
			6256: dout = 12'hfa0;
			6257: dout = 12'hfa0;
			6258: dout = 12'he60;
			6259: dout = 12'h000;
			6260: dout = 12'ha40;
			6261: dout = 12'hfa0;
			6262: dout = 12'hfa0;
			6263: dout = 12'h500;
			6264: dout = 12'h000;
			6265: dout = 12'h000;
			6266: dout = 12'h000;
			6267: dout = 12'h000;
			6268: dout = 12'h000;
			6269: dout = 12'h000;
			6270: dout = 12'h000;
			6271: dout = 12'h000;
			6272: dout = 12'h000;
			6273: dout = 12'h000;
			6274: dout = 12'h000;
			6275: dout = 12'h000;
			6276: dout = 12'h000;
			6277: dout = 12'h000;
			6278: dout = 12'h000;
			6279: dout = 12'h000;
			6280: dout = 12'h000;
			6281: dout = 12'h000;
			6282: dout = 12'h000;
			6283: dout = 12'h000;
			6284: dout = 12'h710;
			6285: dout = 12'hfa0;
			6286: dout = 12'hfa0;
			6287: dout = 12'h930;
			6288: dout = 12'h000;
			6289: dout = 12'h000;
			6290: dout = 12'h000;
			6291: dout = 12'h000;
			6292: dout = 12'h000;
			6293: dout = 12'h000;
			6294: dout = 12'h000;
			6295: dout = 12'h000;
			6296: dout = 12'h000;
			6297: dout = 12'h000;
			6298: dout = 12'h000;
			6299: dout = 12'h400;
			6300: dout = 12'hfa0;
			6301: dout = 12'hfa0;
			6302: dout = 12'hc40;
			6303: dout = 12'h000;
			6304: dout = 12'h000;
			6305: dout = 12'h000;
			6306: dout = 12'h000;
			6307: dout = 12'hd60;
			6308: dout = 12'hfa0;
			6309: dout = 12'hfb0;
			6310: dout = 12'h300;
			6311: dout = 12'h000;
			6312: dout = 12'h000;
			6313: dout = 12'hc50;
			6314: dout = 12'hfa0;
			6315: dout = 12'hfb0;
			6316: dout = 12'h400;
			6317: dout = 12'h000;
			6318: dout = 12'h000;
			6319: dout = 12'h000;
			6320: dout = 12'h200;
			6321: dout = 12'hf90;
			6322: dout = 12'hfa0;
			6323: dout = 12'he60;
			6324: dout = 12'h000;
			6325: dout = 12'h000;
			6326: dout = 12'h000;
			6327: dout = 12'h000;
			6328: dout = 12'h000;
			6329: dout = 12'h000;
			6330: dout = 12'h000;
			6331: dout = 12'h000;
			6332: dout = 12'h000;
			6333: dout = 12'h000;
			6334: dout = 12'h000;
			6335: dout = 12'h000;
			6336: dout = 12'h000;
			6337: dout = 12'h930;
			6338: dout = 12'hfa0;
			6339: dout = 12'hfa0;
			6340: dout = 12'h720;
			6341: dout = 12'h000;
			6342: dout = 12'h000;
			6343: dout = 12'h000;
			6344: dout = 12'h000;
			6345: dout = 12'h000;
			6346: dout = 12'h720;
			6347: dout = 12'hfb0;
			6348: dout = 12'hfb0;
			6349: dout = 12'h930;
			6350: dout = 12'h000;
			6351: dout = 12'h000;
			6352: dout = 12'h000;
			6353: dout = 12'h000;
			6354: dout = 12'h000;
			6355: dout = 12'h000;
			6356: dout = 12'h000;
			6357: dout = 12'h000;

			6358: dout = 12'h000;
			6359: dout = 12'h000;
			6360: dout = 12'h930;
			6361: dout = 12'hfb0;
			6362: dout = 12'hfb0;
			6363: dout = 12'h720;
			6364: dout = 12'h000;
			6365: dout = 12'h000;
			6366: dout = 12'h000;
			6367: dout = 12'h000;
			6368: dout = 12'h000;
			6369: dout = 12'h000;
			6370: dout = 12'h000;
			6371: dout = 12'h000;
			6372: dout = 12'h000;
			6373: dout = 12'h000;
			6374: dout = 12'he80;
			6375: dout = 12'hfb0;
			6376: dout = 12'hfa0;
			6377: dout = 12'h100;
			6378: dout = 12'h610;
			6379: dout = 12'hfb0;
			6380: dout = 12'hfb0;
			6381: dout = 12'ha40;
			6382: dout = 12'h000;
			6383: dout = 12'h000;
			6384: dout = 12'h000;
			6385: dout = 12'h000;
			6386: dout = 12'h000;
			6387: dout = 12'h000;
			6388: dout = 12'h000;
			6389: dout = 12'hd60;
			6390: dout = 12'hfb0;
			6391: dout = 12'hfb0;
			6392: dout = 12'h200;
			6393: dout = 12'h300;
			6394: dout = 12'hfb0;
			6395: dout = 12'hfb0;
			6396: dout = 12'hc50;
			6397: dout = 12'h000;
			6398: dout = 12'h000;
			6399: dout = 12'h000;
			6400: dout = 12'h000;
			6401: dout = 12'h000;
			6402: dout = 12'h000;
			6403: dout = 12'h000;
			6404: dout = 12'h000;
			6405: dout = 12'h200;
			6406: dout = 12'hfb0;
			6407: dout = 12'hfb0;
			6408: dout = 12'he70;
			6409: dout = 12'h000;
			6410: dout = 12'ha40;
			6411: dout = 12'hfb0;
			6412: dout = 12'hfb0;
			6413: dout = 12'h500;
			6414: dout = 12'h000;
			6415: dout = 12'h000;
			6416: dout = 12'h000;
			6417: dout = 12'h000;
			6418: dout = 12'h000;
			6419: dout = 12'h000;
			6420: dout = 12'h000;
			6421: dout = 12'h000;
			6422: dout = 12'h000;
			6423: dout = 12'h000;
			6424: dout = 12'h000;
			6425: dout = 12'h000;
			6426: dout = 12'h000;
			6427: dout = 12'h000;
			6428: dout = 12'h000;
			6429: dout = 12'h000;
			6430: dout = 12'h000;
			6431: dout = 12'h000;
			6432: dout = 12'h000;
			6433: dout = 12'h000;
			6434: dout = 12'h710;
			6435: dout = 12'hfb0;
			6436: dout = 12'hfb0;
			6437: dout = 12'h930;
			6438: dout = 12'h000;
			6439: dout = 12'h000;
			6440: dout = 12'h000;
			6441: dout = 12'h000;
			6442: dout = 12'h000;
			6443: dout = 12'h000;
			6444: dout = 12'h000;
			6445: dout = 12'h000;
			6446: dout = 12'h000;
			6447: dout = 12'h000;
			6448: dout = 12'h000;
			6449: dout = 12'h400;
			6450: dout = 12'hfc0;
			6451: dout = 12'hfb0;
			6452: dout = 12'hc50;
			6453: dout = 12'h000;
			6454: dout = 12'h000;
			6455: dout = 12'h000;
			6456: dout = 12'h000;
			6457: dout = 12'hd50;
			6458: dout = 12'hf80;
			6459: dout = 12'hf90;
			6460: dout = 12'h400;
			6461: dout = 12'h000;
			6462: dout = 12'h000;
			6463: dout = 12'hc40;
			6464: dout = 12'hf80;
			6465: dout = 12'hf90;
			6466: dout = 12'h400;
			6467: dout = 12'h000;
			6468: dout = 12'h000;
			6469: dout = 12'h000;
			6470: dout = 12'h200;
			6471: dout = 12'hfa0;
			6472: dout = 12'hfb0;
			6473: dout = 12'he70;
			6474: dout = 12'h000;
			6475: dout = 12'h000;
			6476: dout = 12'h000;
			6477: dout = 12'h000;
			6478: dout = 12'h000;
			6479: dout = 12'h000;
			6480: dout = 12'h000;
			6481: dout = 12'h000;
			6482: dout = 12'h000;
			6483: dout = 12'h000;
			6484: dout = 12'h000;
			6485: dout = 12'h000;
			6486: dout = 12'h000;
			6487: dout = 12'h930;
			6488: dout = 12'hfb0;
			6489: dout = 12'hfb0;
			6490: dout = 12'h720;
			6491: dout = 12'h000;
			6492: dout = 12'h000;
			6493: dout = 12'h000;
			6494: dout = 12'h000;
			6495: dout = 12'h000;
			6496: dout = 12'h820;
			6497: dout = 12'hf90;
			6498: dout = 12'hf90;
			6499: dout = 12'h920;
			6500: dout = 12'h000;
			6501: dout = 12'h100;
			6502: dout = 12'h100;
			6503: dout = 12'h000;
			6504: dout = 12'h000;
			6505: dout = 12'h000;
			6506: dout = 12'h000;
			6507: dout = 12'h000;

			6508: dout = 12'h000;
			6509: dout = 12'h000;
			6510: dout = 12'h930;
			6511: dout = 12'hfc0;
			6512: dout = 12'hfc0;
			6513: dout = 12'h720;
			6514: dout = 12'h000;
			6515: dout = 12'h000;
			6516: dout = 12'h000;
			6517: dout = 12'h000;
			6518: dout = 12'h000;
			6519: dout = 12'h000;
			6520: dout = 12'h000;
			6521: dout = 12'h000;
			6522: dout = 12'h000;
			6523: dout = 12'h000;
			6524: dout = 12'he80;
			6525: dout = 12'hfc0;
			6526: dout = 12'hfa0;
			6527: dout = 12'h100;
			6528: dout = 12'h610;
			6529: dout = 12'hfc0;
			6530: dout = 12'hfc0;
			6531: dout = 12'ha40;
			6532: dout = 12'h000;
			6533: dout = 12'h000;
			6534: dout = 12'h000;
			6535: dout = 12'h000;
			6536: dout = 12'h000;
			6537: dout = 12'h000;
			6538: dout = 12'h000;
			6539: dout = 12'hd70;
			6540: dout = 12'hfc0;
			6541: dout = 12'hfc0;
			6542: dout = 12'h200;
			6543: dout = 12'h300;
			6544: dout = 12'hfc0;
			6545: dout = 12'hfc0;
			6546: dout = 12'hc60;
			6547: dout = 12'h000;
			6548: dout = 12'h000;
			6549: dout = 12'h000;
			6550: dout = 12'h000;
			6551: dout = 12'h000;
			6552: dout = 12'h000;
			6553: dout = 12'h000;
			6554: dout = 12'h000;
			6555: dout = 12'h200;
			6556: dout = 12'hfc0;
			6557: dout = 12'hfc0;
			6558: dout = 12'he70;
			6559: dout = 12'h000;
			6560: dout = 12'ha40;
			6561: dout = 12'hfc0;
			6562: dout = 12'hfc0;
			6563: dout = 12'h510;
			6564: dout = 12'h000;
			6565: dout = 12'h000;
			6566: dout = 12'h000;
			6567: dout = 12'h000;
			6568: dout = 12'h000;
			6569: dout = 12'h000;
			6570: dout = 12'h000;
			6571: dout = 12'h000;
			6572: dout = 12'h000;
			6573: dout = 12'h000;
			6574: dout = 12'h000;
			6575: dout = 12'h000;
			6576: dout = 12'h000;
			6577: dout = 12'h000;
			6578: dout = 12'h000;
			6579: dout = 12'h000;
			6580: dout = 12'h000;
			6581: dout = 12'h000;
			6582: dout = 12'h000;
			6583: dout = 12'h000;
			6584: dout = 12'h710;
			6585: dout = 12'hfc0;
			6586: dout = 12'hfc0;
			6587: dout = 12'h930;
			6588: dout = 12'h000;
			6589: dout = 12'h000;
			6590: dout = 12'h000;
			6591: dout = 12'h000;
			6592: dout = 12'h000;
			6593: dout = 12'h000;
			6594: dout = 12'h000;
			6595: dout = 12'h000;
			6596: dout = 12'h000;
			6597: dout = 12'h000;
			6598: dout = 12'h000;
			6599: dout = 12'h400;
			6600: dout = 12'hfd0;
			6601: dout = 12'hfc0;
			6602: dout = 12'hc50;
			6603: dout = 12'h000;
			6604: dout = 12'h000;
			6605: dout = 12'h000;
			6606: dout = 12'h000;
			6607: dout = 12'h000;
			6608: dout = 12'h000;
			6609: dout = 12'h000;
			6610: dout = 12'hc50;
			6611: dout = 12'hfa0;
			6612: dout = 12'hfb0;
			6613: dout = 12'h300;
			6614: dout = 12'h000;
			6615: dout = 12'h000;
			6616: dout = 12'h000;
			6617: dout = 12'h000;
			6618: dout = 12'h000;
			6619: dout = 12'h000;
			6620: dout = 12'h200;
			6621: dout = 12'hfb0;
			6622: dout = 12'hfc0;
			6623: dout = 12'he70;
			6624: dout = 12'h000;
			6625: dout = 12'h000;
			6626: dout = 12'h000;
			6627: dout = 12'h000;
			6628: dout = 12'h000;
			6629: dout = 12'h000;
			6630: dout = 12'h000;
			6631: dout = 12'h000;
			6632: dout = 12'h000;
			6633: dout = 12'h000;
			6634: dout = 12'h000;
			6635: dout = 12'h000;
			6636: dout = 12'h000;
			6637: dout = 12'h930;
			6638: dout = 12'hfc0;
			6639: dout = 12'hfc0;
			6640: dout = 12'h720;
			6641: dout = 12'h000;
			6642: dout = 12'h000;
			6643: dout = 12'h000;
			6644: dout = 12'h000;
			6645: dout = 12'h000;
			6646: dout = 12'h000;
			6647: dout = 12'h100;
			6648: dout = 12'h000;
			6649: dout = 12'h710;
			6650: dout = 12'hfa0;
			6651: dout = 12'hfa0;
			6652: dout = 12'ha30;
			6653: dout = 12'h000;
			6654: dout = 12'h000;
			6655: dout = 12'h000;
			6656: dout = 12'h000;
			6657: dout = 12'h000;

			6658: dout = 12'h000;
			6659: dout = 12'h000;
			6660: dout = 12'h940;
			6661: dout = 12'hfe0;
			6662: dout = 12'hfe0;
			6663: dout = 12'h720;
			6664: dout = 12'h000;
			6665: dout = 12'h000;
			6666: dout = 12'h000;
			6667: dout = 12'h000;
			6668: dout = 12'h000;
			6669: dout = 12'h000;
			6670: dout = 12'h000;
			6671: dout = 12'h000;
			6672: dout = 12'h000;
			6673: dout = 12'h000;
			6674: dout = 12'he90;
			6675: dout = 12'hfd0;
			6676: dout = 12'hfc0;
			6677: dout = 12'h100;
			6678: dout = 12'h610;
			6679: dout = 12'hfd0;
			6680: dout = 12'hfd0;
			6681: dout = 12'ha40;
			6682: dout = 12'h000;
			6683: dout = 12'h000;
			6684: dout = 12'h000;
			6685: dout = 12'h000;
			6686: dout = 12'h000;
			6687: dout = 12'h000;
			6688: dout = 12'h000;
			6689: dout = 12'hd70;
			6690: dout = 12'hfd0;
			6691: dout = 12'hfd0;
			6692: dout = 12'h200;
			6693: dout = 12'h300;
			6694: dout = 12'hfd0;
			6695: dout = 12'hfd0;
			6696: dout = 12'hc60;
			6697: dout = 12'h000;
			6698: dout = 12'h000;
			6699: dout = 12'h000;
			6700: dout = 12'h000;
			6701: dout = 12'h000;
			6702: dout = 12'h000;
			6703: dout = 12'h000;
			6704: dout = 12'h000;
			6705: dout = 12'h200;
			6706: dout = 12'hfd0;
			6707: dout = 12'hfd0;
			6708: dout = 12'he80;
			6709: dout = 12'h000;
			6710: dout = 12'ha50;
			6711: dout = 12'hfd0;
			6712: dout = 12'hfd0;
			6713: dout = 12'h510;
			6714: dout = 12'h000;
			6715: dout = 12'h000;
			6716: dout = 12'h000;
			6717: dout = 12'h000;
			6718: dout = 12'h000;
			6719: dout = 12'h000;
			6720: dout = 12'h000;
			6721: dout = 12'h000;
			6722: dout = 12'h000;
			6723: dout = 12'h000;
			6724: dout = 12'h000;
			6725: dout = 12'h000;
			6726: dout = 12'h000;
			6727: dout = 12'h000;
			6728: dout = 12'h000;
			6729: dout = 12'h000;
			6730: dout = 12'h000;
			6731: dout = 12'h000;
			6732: dout = 12'h000;
			6733: dout = 12'h000;
			6734: dout = 12'h720;
			6735: dout = 12'hfe0;
			6736: dout = 12'hfe0;
			6737: dout = 12'h940;
			6738: dout = 12'h000;
			6739: dout = 12'h000;
			6740: dout = 12'h000;
			6741: dout = 12'h000;
			6742: dout = 12'h000;
			6743: dout = 12'h000;
			6744: dout = 12'h000;
			6745: dout = 12'h000;
			6746: dout = 12'h000;
			6747: dout = 12'h000;
			6748: dout = 12'h000;
			6749: dout = 12'h400;
			6750: dout = 12'hfe0;
			6751: dout = 12'hfe0;
			6752: dout = 12'hc60;
			6753: dout = 12'h000;
			6754: dout = 12'h000;
			6755: dout = 12'h000;
			6756: dout = 12'h000;
			6757: dout = 12'h000;
			6758: dout = 12'h000;
			6759: dout = 12'h000;
			6760: dout = 12'hd70;
			6761: dout = 12'hfd0;
			6762: dout = 12'hfe0;
			6763: dout = 12'h300;
			6764: dout = 12'h000;
			6765: dout = 12'h000;
			6766: dout = 12'h000;
			6767: dout = 12'h000;
			6768: dout = 12'h000;
			6769: dout = 12'h000;
			6770: dout = 12'h200;
			6771: dout = 12'hfc0;
			6772: dout = 12'hfd0;
			6773: dout = 12'he80;
			6774: dout = 12'h000;
			6775: dout = 12'h000;
			6776: dout = 12'h000;
			6777: dout = 12'h000;
			6778: dout = 12'h000;
			6779: dout = 12'h000;
			6780: dout = 12'h000;
			6781: dout = 12'h000;
			6782: dout = 12'h000;
			6783: dout = 12'h000;
			6784: dout = 12'h000;
			6785: dout = 12'h000;
			6786: dout = 12'h000;
			6787: dout = 12'h930;
			6788: dout = 12'hfd0;
			6789: dout = 12'hfd0;
			6790: dout = 12'h720;
			6791: dout = 12'h000;
			6792: dout = 12'h000;
			6793: dout = 12'h000;
			6794: dout = 12'h000;
			6795: dout = 12'h000;
			6796: dout = 12'h000;
			6797: dout = 12'h000;
			6798: dout = 12'h000;
			6799: dout = 12'h720;
			6800: dout = 12'hfe0;
			6801: dout = 12'hfe0;
			6802: dout = 12'h940;
			6803: dout = 12'h000;
			6804: dout = 12'h000;
			6805: dout = 12'h000;
			6806: dout = 12'h000;
			6807: dout = 12'h000;

			6808: dout = 12'h000;
			6809: dout = 12'h000;
			6810: dout = 12'h930;
			6811: dout = 12'hfa0;
			6812: dout = 12'hfa0;
			6813: dout = 12'h710;
			6814: dout = 12'h100;
			6815: dout = 12'h200;
			6816: dout = 12'h200;
			6817: dout = 12'h200;
			6818: dout = 12'h200;
			6819: dout = 12'h200;
			6820: dout = 12'h200;
			6821: dout = 12'h200;
			6822: dout = 12'h100;
			6823: dout = 12'h200;
			6824: dout = 12'hd70;
			6825: dout = 12'hea0;
			6826: dout = 12'he90;
			6827: dout = 12'h100;
			6828: dout = 12'h610;
			6829: dout = 12'hfe0;
			6830: dout = 12'hfe0;
			6831: dout = 12'ha50;
			6832: dout = 12'h000;
			6833: dout = 12'h000;
			6834: dout = 12'h000;
			6835: dout = 12'h000;
			6836: dout = 12'h000;
			6837: dout = 12'h000;
			6838: dout = 12'h000;
			6839: dout = 12'hd80;
			6840: dout = 12'hfe0;
			6841: dout = 12'hfe0;
			6842: dout = 12'h200;
			6843: dout = 12'h300;
			6844: dout = 12'hfe0;
			6845: dout = 12'hfe0;
			6846: dout = 12'hc70;
			6847: dout = 12'h000;
			6848: dout = 12'h000;
			6849: dout = 12'h000;
			6850: dout = 12'h000;
			6851: dout = 12'h000;
			6852: dout = 12'h000;
			6853: dout = 12'h000;
			6854: dout = 12'h000;
			6855: dout = 12'h200;
			6856: dout = 12'hfe0;
			6857: dout = 12'hfe0;
			6858: dout = 12'he80;
			6859: dout = 12'h000;
			6860: dout = 12'ha50;
			6861: dout = 12'hfe0;
			6862: dout = 12'hff0;
			6863: dout = 12'h600;
			6864: dout = 12'h100;
			6865: dout = 12'h200;
			6866: dout = 12'h200;
			6867: dout = 12'h200;
			6868: dout = 12'h200;
			6869: dout = 12'h200;
			6870: dout = 12'h200;
			6871: dout = 12'h200;
			6872: dout = 12'h200;
			6873: dout = 12'h200;
			6874: dout = 12'h200;
			6875: dout = 12'h100;
			6876: dout = 12'h000;
			6877: dout = 12'h000;
			6878: dout = 12'h000;
			6879: dout = 12'h000;
			6880: dout = 12'h000;
			6881: dout = 12'h000;
			6882: dout = 12'h000;
			6883: dout = 12'h000;
			6884: dout = 12'h710;
			6885: dout = 12'hfa0;
			6886: dout = 12'hea0;
			6887: dout = 12'h930;
			6888: dout = 12'h100;
			6889: dout = 12'h200;
			6890: dout = 12'h200;
			6891: dout = 12'h200;
			6892: dout = 12'h200;
			6893: dout = 12'h200;
			6894: dout = 12'h200;
			6895: dout = 12'h200;
			6896: dout = 12'h200;
			6897: dout = 12'h200;
			6898: dout = 12'h100;
			6899: dout = 12'h500;
			6900: dout = 12'hfa0;
			6901: dout = 12'hea0;
			6902: dout = 12'hc40;
			6903: dout = 12'h000;
			6904: dout = 12'h000;
			6905: dout = 12'h000;
			6906: dout = 12'h000;
			6907: dout = 12'h000;
			6908: dout = 12'h000;
			6909: dout = 12'h000;
			6910: dout = 12'hd70;
			6911: dout = 12'hfe0;
			6912: dout = 12'hff0;
			6913: dout = 12'h300;
			6914: dout = 12'h000;
			6915: dout = 12'h000;
			6916: dout = 12'h000;
			6917: dout = 12'h000;
			6918: dout = 12'h000;
			6919: dout = 12'h000;
			6920: dout = 12'h200;
			6921: dout = 12'hfd0;
			6922: dout = 12'hfe0;
			6923: dout = 12'hd80;
			6924: dout = 12'h100;
			6925: dout = 12'h100;
			6926: dout = 12'h200;
			6927: dout = 12'h200;
			6928: dout = 12'h200;
			6929: dout = 12'h200;
			6930: dout = 12'h200;
			6931: dout = 12'h200;
			6932: dout = 12'h200;
			6933: dout = 12'h200;
			6934: dout = 12'h200;
			6935: dout = 12'h200;
			6936: dout = 12'h000;
			6937: dout = 12'h940;
			6938: dout = 12'hfe0;
			6939: dout = 12'hfe0;
			6940: dout = 12'h730;
			6941: dout = 12'h000;
			6942: dout = 12'h000;
			6943: dout = 12'h000;
			6944: dout = 12'h000;
			6945: dout = 12'h000;
			6946: dout = 12'h000;
			6947: dout = 12'h000;
			6948: dout = 12'h000;
			6949: dout = 12'h720;
			6950: dout = 12'hfa0;
			6951: dout = 12'hea0;
			6952: dout = 12'h930;
			6953: dout = 12'h100;
			6954: dout = 12'h200;
			6955: dout = 12'h200;
			6956: dout = 12'h000;
			6957: dout = 12'h000;

			6958: dout = 12'h000;
			6959: dout = 12'h000;
			6960: dout = 12'h000;
			6961: dout = 12'h000;
			6962: dout = 12'h000;
			6963: dout = 12'h830;
			6964: dout = 12'hfe0;
			6965: dout = 12'hfd0;
			6966: dout = 12'hfd0;
			6967: dout = 12'hfd0;
			6968: dout = 12'hfd0;
			6969: dout = 12'hfd0;
			6970: dout = 12'hfd0;
			6971: dout = 12'hfd0;
			6972: dout = 12'hfd0;
			6973: dout = 12'hfc0;
			6974: dout = 12'h100;
			6975: dout = 12'h000;
			6976: dout = 12'h000;
			6977: dout = 12'h000;
			6978: dout = 12'h610;
			6979: dout = 12'hff0;
			6980: dout = 12'hff0;
			6981: dout = 12'ha50;
			6982: dout = 12'h000;
			6983: dout = 12'h000;
			6984: dout = 12'h000;
			6985: dout = 12'h000;
			6986: dout = 12'h000;
			6987: dout = 12'h000;
			6988: dout = 12'h000;
			6989: dout = 12'hd80;
			6990: dout = 12'hff0;
			6991: dout = 12'hff0;
			6992: dout = 12'h200;
			6993: dout = 12'h300;
			6994: dout = 12'hff0;
			6995: dout = 12'hff0;
			6996: dout = 12'hc70;
			6997: dout = 12'h000;
			6998: dout = 12'h000;
			6999: dout = 12'h000;
			7000: dout = 12'h000;
			7001: dout = 12'h000;
			7002: dout = 12'h000;
			7003: dout = 12'h000;
			7004: dout = 12'h000;
			7005: dout = 12'h200;
			7006: dout = 12'hff0;
			7007: dout = 12'hff0;
			7008: dout = 12'he90;
			7009: dout = 12'h000;
			7010: dout = 12'ha50;
			7011: dout = 12'hff0;
			7012: dout = 12'hfe0;
			7013: dout = 12'hfd0;
			7014: dout = 12'hfd0;
			7015: dout = 12'hfd0;
			7016: dout = 12'hfd0;
			7017: dout = 12'hfd0;
			7018: dout = 12'hfd0;
			7019: dout = 12'hfd0;
			7020: dout = 12'hfd0;
			7021: dout = 12'hfd0;
			7022: dout = 12'hfd0;
			7023: dout = 12'hfd0;
			7024: dout = 12'hfe0;
			7025: dout = 12'h820;
			7026: dout = 12'h000;
			7027: dout = 12'h000;
			7028: dout = 12'h000;
			7029: dout = 12'h000;
			7030: dout = 12'h000;
			7031: dout = 12'h000;
			7032: dout = 12'h000;
			7033: dout = 12'h000;
			7034: dout = 12'h000;
			7035: dout = 12'h000;
			7036: dout = 12'h000;
			7037: dout = 12'h610;
			7038: dout = 12'hfe0;
			7039: dout = 12'hfd0;
			7040: dout = 12'hfd0;
			7041: dout = 12'hfd0;
			7042: dout = 12'hfd0;
			7043: dout = 12'hfd0;
			7044: dout = 12'hfd0;
			7045: dout = 12'hfd0;
			7046: dout = 12'hfd0;
			7047: dout = 12'hfd0;
			7048: dout = 12'hfe0;
			7049: dout = 12'hb60;
			7050: dout = 12'h000;
			7051: dout = 12'h000;
			7052: dout = 12'h000;
			7053: dout = 12'h000;
			7054: dout = 12'h000;
			7055: dout = 12'h000;
			7056: dout = 12'h000;
			7057: dout = 12'h000;
			7058: dout = 12'h000;
			7059: dout = 12'h000;
			7060: dout = 12'hd80;
			7061: dout = 12'hff0;
			7062: dout = 12'hff0;
			7063: dout = 12'h300;
			7064: dout = 12'h000;
			7065: dout = 12'h000;
			7066: dout = 12'h000;
			7067: dout = 12'h000;
			7068: dout = 12'h000;
			7069: dout = 12'h000;
			7070: dout = 12'h200;
			7071: dout = 12'hfe0;
			7072: dout = 12'hfe0;
			7073: dout = 12'hfe0;
			7074: dout = 12'hfd0;
			7075: dout = 12'hfd0;
			7076: dout = 12'hfd0;
			7077: dout = 12'hfd0;
			7078: dout = 12'hfd0;
			7079: dout = 12'hfd0;
			7080: dout = 12'hfd0;
			7081: dout = 12'hfd0;
			7082: dout = 12'hfd0;
			7083: dout = 12'hfd0;
			7084: dout = 12'hfe0;
			7085: dout = 12'hfa0;
			7086: dout = 12'h000;
			7087: dout = 12'h840;
			7088: dout = 12'hff0;
			7089: dout = 12'hff0;
			7090: dout = 12'h730;
			7091: dout = 12'h000;
			7092: dout = 12'h000;
			7093: dout = 12'h000;
			7094: dout = 12'h000;
			7095: dout = 12'h000;
			7096: dout = 12'h000;
			7097: dout = 12'h000;
			7098: dout = 12'h000;
			7099: dout = 12'h000;
			7100: dout = 12'h000;
			7101: dout = 12'h000;
			7102: dout = 12'h610;
			7103: dout = 12'hfe0;
			7104: dout = 12'hfe0;
			7105: dout = 12'ha50;
			7106: dout = 12'h000;
			7107: dout = 12'h000;

			7108: dout = 12'h000;
			7109: dout = 12'h000;
			7110: dout = 12'h000;
			7111: dout = 12'h000;
			7112: dout = 12'h000;
			7113: dout = 12'h940;
			7114: dout = 12'hff0;
			7115: dout = 12'hff0;
			7116: dout = 12'hff0;
			7117: dout = 12'hff0;
			7118: dout = 12'hff0;
			7119: dout = 12'hff0;
			7120: dout = 12'hff0;
			7121: dout = 12'hff0;
			7122: dout = 12'hff0;
			7123: dout = 12'hfe0;
			7124: dout = 12'h100;
			7125: dout = 12'h000;
			7126: dout = 12'h000;
			7127: dout = 12'h000;
			7128: dout = 12'h620;
			7129: dout = 12'hff0;
			7130: dout = 12'hff0;
			7131: dout = 12'ha60;
			7132: dout = 12'h000;
			7133: dout = 12'h000;
			7134: dout = 12'h000;
			7135: dout = 12'h000;
			7136: dout = 12'h000;
			7137: dout = 12'h000;
			7138: dout = 12'h000;
			7139: dout = 12'hd90;
			7140: dout = 12'hff0;
			7141: dout = 12'hff0;
			7142: dout = 12'h200;
			7143: dout = 12'h300;
			7144: dout = 12'hff0;
			7145: dout = 12'hff0;
			7146: dout = 12'hc80;
			7147: dout = 12'h000;
			7148: dout = 12'h000;
			7149: dout = 12'h000;
			7150: dout = 12'h000;
			7151: dout = 12'h000;
			7152: dout = 12'h000;
			7153: dout = 12'h000;
			7154: dout = 12'h000;
			7155: dout = 12'h200;
			7156: dout = 12'hff0;
			7157: dout = 12'hff0;
			7158: dout = 12'hea0;
			7159: dout = 12'h000;
			7160: dout = 12'hb60;
			7161: dout = 12'hff0;
			7162: dout = 12'hff0;
			7163: dout = 12'hff0;
			7164: dout = 12'hff0;
			7165: dout = 12'hff0;
			7166: dout = 12'hff0;
			7167: dout = 12'hff0;
			7168: dout = 12'hff0;
			7169: dout = 12'hff0;
			7170: dout = 12'hff0;
			7171: dout = 12'hff0;
			7172: dout = 12'hff0;
			7173: dout = 12'hff0;
			7174: dout = 12'hff0;
			7175: dout = 12'h830;
			7176: dout = 12'h000;
			7177: dout = 12'h000;
			7178: dout = 12'h000;
			7179: dout = 12'h000;
			7180: dout = 12'h000;
			7181: dout = 12'h000;
			7182: dout = 12'h000;
			7183: dout = 12'h000;
			7184: dout = 12'h000;
			7185: dout = 12'h000;
			7186: dout = 12'h000;
			7187: dout = 12'h610;
			7188: dout = 12'hff0;
			7189: dout = 12'hff0;
			7190: dout = 12'hff0;
			7191: dout = 12'hff0;
			7192: dout = 12'hff0;
			7193: dout = 12'hff0;
			7194: dout = 12'hff0;
			7195: dout = 12'hff0;
			7196: dout = 12'hff0;
			7197: dout = 12'hff0;
			7198: dout = 12'hff0;
			7199: dout = 12'hb70;
			7200: dout = 12'h000;
			7201: dout = 12'h000;
			7202: dout = 12'h000;
			7203: dout = 12'h000;
			7204: dout = 12'h000;
			7205: dout = 12'h000;
			7206: dout = 12'h000;
			7207: dout = 12'h000;
			7208: dout = 12'h000;
			7209: dout = 12'h000;
			7210: dout = 12'hd90;
			7211: dout = 12'hff0;
			7212: dout = 12'hff0;
			7213: dout = 12'h300;
			7214: dout = 12'h000;
			7215: dout = 12'h000;
			7216: dout = 12'h000;
			7217: dout = 12'h000;
			7218: dout = 12'h000;
			7219: dout = 12'h000;
			7220: dout = 12'h200;
			7221: dout = 12'hff0;
			7222: dout = 12'hff0;
			7223: dout = 12'hff0;
			7224: dout = 12'hff0;
			7225: dout = 12'hff0;
			7226: dout = 12'hff0;
			7227: dout = 12'hff0;
			7228: dout = 12'hff0;
			7229: dout = 12'hff0;
			7230: dout = 12'hff0;
			7231: dout = 12'hff0;
			7232: dout = 12'hff0;
			7233: dout = 12'hff0;
			7234: dout = 12'hff0;
			7235: dout = 12'hfc0;
			7236: dout = 12'h000;
			7237: dout = 12'h840;
			7238: dout = 12'hff0;
			7239: dout = 12'hff0;
			7240: dout = 12'h830;
			7241: dout = 12'h000;
			7242: dout = 12'h000;
			7243: dout = 12'h000;
			7244: dout = 12'h000;
			7245: dout = 12'h000;
			7246: dout = 12'h000;
			7247: dout = 12'h000;
			7248: dout = 12'h000;
			7249: dout = 12'h000;
			7250: dout = 12'h000;
			7251: dout = 12'h000;
			7252: dout = 12'h620;
			7253: dout = 12'hff0;
			7254: dout = 12'hff0;
			7255: dout = 12'ha60;
			7256: dout = 12'h000;
			7257: dout = 12'h000;

			7258: dout = 12'h000;
			7259: dout = 12'h000;
			7260: dout = 12'h000;
			7261: dout = 12'h000;
			7262: dout = 12'h000;
			7263: dout = 12'h830;
			7264: dout = 12'hea0;
			7265: dout = 12'hda0;
			7266: dout = 12'hda0;
			7267: dout = 12'hda0;
			7268: dout = 12'hda0;
			7269: dout = 12'hda0;
			7270: dout = 12'hda0;
			7271: dout = 12'hda0;
			7272: dout = 12'hda0;
			7273: dout = 12'he90;
			7274: dout = 12'h200;
			7275: dout = 12'h000;
			7276: dout = 12'h000;
			7277: dout = 12'h000;
			7278: dout = 12'h610;
			7279: dout = 12'hea0;
			7280: dout = 12'hea0;
			7281: dout = 12'ha40;
			7282: dout = 12'h000;
			7283: dout = 12'h000;
			7284: dout = 12'h000;
			7285: dout = 12'h000;
			7286: dout = 12'h000;
			7287: dout = 12'h000;
			7288: dout = 12'h000;
			7289: dout = 12'hc60;
			7290: dout = 12'hea0;
			7291: dout = 12'hea0;
			7292: dout = 12'h300;
			7293: dout = 12'h400;
			7294: dout = 12'hea0;
			7295: dout = 12'hea0;
			7296: dout = 12'hb50;
			7297: dout = 12'h000;
			7298: dout = 12'h000;
			7299: dout = 12'h000;
			7300: dout = 12'h000;
			7301: dout = 12'h000;
			7302: dout = 12'h000;
			7303: dout = 12'h000;
			7304: dout = 12'h000;
			7305: dout = 12'h300;
			7306: dout = 12'hea0;
			7307: dout = 12'hea0;
			7308: dout = 12'hd60;
			7309: dout = 12'h000;
			7310: dout = 12'ha40;
			7311: dout = 12'hea0;
			7312: dout = 12'hda0;
			7313: dout = 12'hda0;
			7314: dout = 12'hda0;
			7315: dout = 12'hda0;
			7316: dout = 12'hda0;
			7317: dout = 12'hda0;
			7318: dout = 12'hda0;
			7319: dout = 12'hda0;
			7320: dout = 12'hda0;
			7321: dout = 12'hda0;
			7322: dout = 12'hda0;
			7323: dout = 12'hda0;
			7324: dout = 12'hea0;
			7325: dout = 12'h820;
			7326: dout = 12'h000;
			7327: dout = 12'h000;
			7328: dout = 12'h000;
			7329: dout = 12'h000;
			7330: dout = 12'h000;
			7331: dout = 12'h000;
			7332: dout = 12'h000;
			7333: dout = 12'h000;
			7334: dout = 12'h000;
			7335: dout = 12'h000;
			7336: dout = 12'h000;
			7337: dout = 12'h710;
			7338: dout = 12'hea0;
			7339: dout = 12'hda0;
			7340: dout = 12'hda0;
			7341: dout = 12'hda0;
			7342: dout = 12'hda0;
			7343: dout = 12'hda0;
			7344: dout = 12'hda0;
			7345: dout = 12'hda0;
			7346: dout = 12'hda0;
			7347: dout = 12'hda0;
			7348: dout = 12'hea0;
			7349: dout = 12'hb40;
			7350: dout = 12'h000;
			7351: dout = 12'h000;
			7352: dout = 12'h000;
			7353: dout = 12'h000;
			7354: dout = 12'h000;
			7355: dout = 12'h000;
			7356: dout = 12'h000;
			7357: dout = 12'h000;
			7358: dout = 12'h000;
			7359: dout = 12'h000;
			7360: dout = 12'hc50;
			7361: dout = 12'hea0;
			7362: dout = 12'heb0;
			7363: dout = 12'h400;
			7364: dout = 12'h000;
			7365: dout = 12'h000;
			7366: dout = 12'h000;
			7367: dout = 12'h000;
			7368: dout = 12'h000;
			7369: dout = 12'h000;
			7370: dout = 12'h300;
			7371: dout = 12'hea0;
			7372: dout = 12'hda0;
			7373: dout = 12'hda0;
			7374: dout = 12'hda0;
			7375: dout = 12'hda0;
			7376: dout = 12'hda0;
			7377: dout = 12'hda0;
			7378: dout = 12'hda0;
			7379: dout = 12'hda0;
			7380: dout = 12'hda0;
			7381: dout = 12'hda0;
			7382: dout = 12'hda0;
			7383: dout = 12'hda0;
			7384: dout = 12'hea0;
			7385: dout = 12'hd80;
			7386: dout = 12'h000;
			7387: dout = 12'h830;
			7388: dout = 12'hea0;
			7389: dout = 12'hea0;
			7390: dout = 12'h820;
			7391: dout = 12'h000;
			7392: dout = 12'h000;
			7393: dout = 12'h000;
			7394: dout = 12'h000;
			7395: dout = 12'h000;
			7396: dout = 12'h000;
			7397: dout = 12'h000;
			7398: dout = 12'h000;
			7399: dout = 12'h000;
			7400: dout = 12'h000;
			7401: dout = 12'h000;
			7402: dout = 12'h610;
			7403: dout = 12'hea0;
			7404: dout = 12'hea0;
			7405: dout = 12'ha30;
			7406: dout = 12'h000;
			7407: dout = 12'h000;

			7408: dout = 12'h000;
			7409: dout = 12'h000;
			7410: dout = 12'h000;
			7411: dout = 12'h000;
			7412: dout = 12'h000;
			7413: dout = 12'h000;
			7414: dout = 12'h000;
			7415: dout = 12'h000;
			7416: dout = 12'h000;
			7417: dout = 12'h000;
			7418: dout = 12'h000;
			7419: dout = 12'h000;
			7420: dout = 12'h000;
			7421: dout = 12'h000;
			7422: dout = 12'h000;
			7423: dout = 12'h000;
			7424: dout = 12'h000;
			7425: dout = 12'h000;
			7426: dout = 12'h000;
			7427: dout = 12'h000;
			7428: dout = 12'h000;
			7429: dout = 12'h000;
			7430: dout = 12'h000;
			7431: dout = 12'h000;
			7432: dout = 12'h000;
			7433: dout = 12'h000;
			7434: dout = 12'h000;
			7435: dout = 12'h000;
			7436: dout = 12'h000;
			7437: dout = 12'h000;
			7438: dout = 12'h000;
			7439: dout = 12'h000;
			7440: dout = 12'h000;
			7441: dout = 12'h000;
			7442: dout = 12'h000;
			7443: dout = 12'h000;
			7444: dout = 12'h000;
			7445: dout = 12'h000;
			7446: dout = 12'h000;
			7447: dout = 12'h000;
			7448: dout = 12'h000;
			7449: dout = 12'h000;
			7450: dout = 12'h000;
			7451: dout = 12'h000;
			7452: dout = 12'h000;
			7453: dout = 12'h000;
			7454: dout = 12'h000;
			7455: dout = 12'h000;
			7456: dout = 12'h000;
			7457: dout = 12'h000;
			7458: dout = 12'h000;
			7459: dout = 12'h000;
			7460: dout = 12'h000;
			7461: dout = 12'h000;
			7462: dout = 12'h000;
			7463: dout = 12'h000;
			7464: dout = 12'h000;
			7465: dout = 12'h000;
			7466: dout = 12'h000;
			7467: dout = 12'h000;
			7468: dout = 12'h000;
			7469: dout = 12'h000;
			7470: dout = 12'h000;
			7471: dout = 12'h000;
			7472: dout = 12'h000;
			7473: dout = 12'h000;
			7474: dout = 12'h000;
			7475: dout = 12'h000;
			7476: dout = 12'h000;
			7477: dout = 12'h000;
			7478: dout = 12'h000;
			7479: dout = 12'h000;
			7480: dout = 12'h000;
			7481: dout = 12'h000;
			7482: dout = 12'h000;
			7483: dout = 12'h000;
			7484: dout = 12'h000;
			7485: dout = 12'h000;
			7486: dout = 12'h000;
			7487: dout = 12'h000;
			7488: dout = 12'h000;
			7489: dout = 12'h000;
			7490: dout = 12'h000;
			7491: dout = 12'h000;
			7492: dout = 12'h000;
			7493: dout = 12'h000;
			7494: dout = 12'h000;
			7495: dout = 12'h000;
			7496: dout = 12'h000;
			7497: dout = 12'h000;
			7498: dout = 12'h000;
			7499: dout = 12'h000;
			7500: dout = 12'h000;
			7501: dout = 12'h000;
			7502: dout = 12'h000;
			7503: dout = 12'h000;
			7504: dout = 12'h000;
			7505: dout = 12'h000;
			7506: dout = 12'h000;
			7507: dout = 12'h000;
			7508: dout = 12'h000;
			7509: dout = 12'h000;
			7510: dout = 12'h000;
			7511: dout = 12'h000;
			7512: dout = 12'h000;
			7513: dout = 12'h000;
			7514: dout = 12'h000;
			7515: dout = 12'h000;
			7516: dout = 12'h000;
			7517: dout = 12'h000;
			7518: dout = 12'h000;
			7519: dout = 12'h000;
			7520: dout = 12'h000;
			7521: dout = 12'h000;
			7522: dout = 12'h000;
			7523: dout = 12'h000;
			7524: dout = 12'h000;
			7525: dout = 12'h000;
			7526: dout = 12'h000;
			7527: dout = 12'h000;
			7528: dout = 12'h000;
			7529: dout = 12'h000;
			7530: dout = 12'h000;
			7531: dout = 12'h000;
			7532: dout = 12'h000;
			7533: dout = 12'h000;
			7534: dout = 12'h000;
			7535: dout = 12'h000;
			7536: dout = 12'h000;
			7537: dout = 12'h000;
			7538: dout = 12'h000;
			7539: dout = 12'h000;
			7540: dout = 12'h000;
			7541: dout = 12'h000;
			7542: dout = 12'h000;
			7543: dout = 12'h000;
			7544: dout = 12'h000;
			7545: dout = 12'h000;
			7546: dout = 12'h000;
			7547: dout = 12'h000;
			7548: dout = 12'h000;
			7549: dout = 12'h000;
			7550: dout = 12'h000;
			7551: dout = 12'h000;
			7552: dout = 12'h000;
			7553: dout = 12'h000;
			7554: dout = 12'h000;
			7555: dout = 12'h000;
			7556: dout = 12'h000;
			7557: dout = 12'h000;

			7558: dout = 12'h000;
			7559: dout = 12'h000;
			7560: dout = 12'h000;
			7561: dout = 12'h000;
			7562: dout = 12'h000;
			7563: dout = 12'h000;
			7564: dout = 12'h000;
			7565: dout = 12'h000;
			7566: dout = 12'h000;
			7567: dout = 12'h000;
			7568: dout = 12'h000;
			7569: dout = 12'h000;
			7570: dout = 12'h000;
			7571: dout = 12'h000;
			7572: dout = 12'h000;
			7573: dout = 12'h000;
			7574: dout = 12'h000;
			7575: dout = 12'h000;
			7576: dout = 12'h000;
			7577: dout = 12'h000;
			7578: dout = 12'h000;
			7579: dout = 12'h000;
			7580: dout = 12'h000;
			7581: dout = 12'h000;
			7582: dout = 12'h000;
			7583: dout = 12'h000;
			7584: dout = 12'h000;
			7585: dout = 12'h000;
			7586: dout = 12'h000;
			7587: dout = 12'h000;
			7588: dout = 12'h000;
			7589: dout = 12'h000;
			7590: dout = 12'h000;
			7591: dout = 12'h000;
			7592: dout = 12'h000;
			7593: dout = 12'h000;
			7594: dout = 12'h000;
			7595: dout = 12'h000;
			7596: dout = 12'h000;
			7597: dout = 12'h000;
			7598: dout = 12'h000;
			7599: dout = 12'h000;
			7600: dout = 12'h000;
			7601: dout = 12'h000;
			7602: dout = 12'h000;
			7603: dout = 12'h000;
			7604: dout = 12'h000;
			7605: dout = 12'h000;
			7606: dout = 12'h000;
			7607: dout = 12'h000;
			7608: dout = 12'h000;
			7609: dout = 12'h000;
			7610: dout = 12'h000;
			7611: dout = 12'h000;
			7612: dout = 12'h000;
			7613: dout = 12'h000;
			7614: dout = 12'h000;
			7615: dout = 12'h000;
			7616: dout = 12'h000;
			7617: dout = 12'h000;
			7618: dout = 12'h000;
			7619: dout = 12'h000;
			7620: dout = 12'h000;
			7621: dout = 12'h000;
			7622: dout = 12'h000;
			7623: dout = 12'h000;
			7624: dout = 12'h000;
			7625: dout = 12'h000;
			7626: dout = 12'h000;
			7627: dout = 12'h000;
			7628: dout = 12'h000;
			7629: dout = 12'h000;
			7630: dout = 12'h000;
			7631: dout = 12'h000;
			7632: dout = 12'h000;
			7633: dout = 12'h000;
			7634: dout = 12'h000;
			7635: dout = 12'h000;
			7636: dout = 12'h000;
			7637: dout = 12'h000;
			7638: dout = 12'h000;
			7639: dout = 12'h000;
			7640: dout = 12'h000;
			7641: dout = 12'h000;
			7642: dout = 12'h000;
			7643: dout = 12'h000;
			7644: dout = 12'h000;
			7645: dout = 12'h000;
			7646: dout = 12'h000;
			7647: dout = 12'h000;
			7648: dout = 12'h000;
			7649: dout = 12'h000;
			7650: dout = 12'h000;
			7651: dout = 12'h000;
			7652: dout = 12'h000;
			7653: dout = 12'h000;
			7654: dout = 12'h000;
			7655: dout = 12'h000;
			7656: dout = 12'h000;
			7657: dout = 12'h000;
			7658: dout = 12'h000;
			7659: dout = 12'h000;
			7660: dout = 12'h000;
			7661: dout = 12'h000;
			7662: dout = 12'h000;
			7663: dout = 12'h000;
			7664: dout = 12'h000;
			7665: dout = 12'h000;
			7666: dout = 12'h000;
			7667: dout = 12'h000;
			7668: dout = 12'h000;
			7669: dout = 12'h000;
			7670: dout = 12'h000;
			7671: dout = 12'h000;
			7672: dout = 12'h000;
			7673: dout = 12'h000;
			7674: dout = 12'h000;
			7675: dout = 12'h000;
			7676: dout = 12'h000;
			7677: dout = 12'h000;
			7678: dout = 12'h000;
			7679: dout = 12'h000;
			7680: dout = 12'h000;
			7681: dout = 12'h000;
			7682: dout = 12'h000;
			7683: dout = 12'h000;
			7684: dout = 12'h000;
			7685: dout = 12'h000;
			7686: dout = 12'h000;
			7687: dout = 12'h000;
			7688: dout = 12'h000;
			7689: dout = 12'h000;
			7690: dout = 12'h000;
			7691: dout = 12'h000;
			7692: dout = 12'h000;
			7693: dout = 12'h000;
			7694: dout = 12'h000;
			7695: dout = 12'h000;
			7696: dout = 12'h000;
			7697: dout = 12'h000;
			7698: dout = 12'h000;
			7699: dout = 12'h000;
			7700: dout = 12'h000;
			7701: dout = 12'h000;
			7702: dout = 12'h000;
			7703: dout = 12'h000;
			7704: dout = 12'h000;
			7705: dout = 12'h000;
			7706: dout = 12'h000;
			7707: dout = 12'h000;

			7708: dout = 12'h000;
			7709: dout = 12'h000;
			7710: dout = 12'h000;
			7711: dout = 12'h000;
			7712: dout = 12'h000;
			7713: dout = 12'h000;
			7714: dout = 12'h000;
			7715: dout = 12'h000;
			7716: dout = 12'h000;
			7717: dout = 12'h110;
			7718: dout = 12'h660;
			7719: dout = 12'h110;
			7720: dout = 12'h000;
			7721: dout = 12'h000;
			7722: dout = 12'h000;
			7723: dout = 12'h000;

			7724: dout = 12'h000;
			7725: dout = 12'h000;
			7726: dout = 12'h000;
			7727: dout = 12'h000;
			7728: dout = 12'h000;
			7729: dout = 12'h000;
			7730: dout = 12'h000;
			7731: dout = 12'h000;
			7732: dout = 12'h000;
			7733: dout = 12'h340;
			7734: dout = 12'hff0;
			7735: dout = 12'h330;
			7736: dout = 12'h000;
			7737: dout = 12'h000;
			7738: dout = 12'h000;
			7739: dout = 12'h000;

			7740: dout = 12'h000;
			7741: dout = 12'h000;
			7742: dout = 12'h000;
			7743: dout = 12'h000;
			7744: dout = 12'h000;
			7745: dout = 12'h000;
			7746: dout = 12'h220;
			7747: dout = 12'hdd0;
			7748: dout = 12'h340;
			7749: dout = 12'h000;
			7750: dout = 12'h220;
			7751: dout = 12'h000;
			7752: dout = 12'h440;
			7753: dout = 12'hdd0;
			7754: dout = 12'h110;
			7755: dout = 12'h000;

			7756: dout = 12'h000;
			7757: dout = 12'h000;
			7758: dout = 12'h000;
			7759: dout = 12'h000;
			7760: dout = 12'h000;
			7761: dout = 12'h000;
			7762: dout = 12'h110;
			7763: dout = 12'haa0;
			7764: dout = 12'h660;
			7765: dout = 12'h540;
			7766: dout = 12'h500;
			7767: dout = 12'h540;
			7768: dout = 12'h670;
			7769: dout = 12'haa0;
			7770: dout = 12'h110;
			7771: dout = 12'h000;

			7772: dout = 12'h000;
			7773: dout = 12'h000;
			7774: dout = 12'h000;
			7775: dout = 12'h000;
			7776: dout = 12'h000;
			7777: dout = 12'h000;
			7778: dout = 12'h000;
			7779: dout = 12'h000;
			7780: dout = 12'hab0;
			7781: dout = 12'hfc0;
			7782: dout = 12'hf00;
			7783: dout = 12'hfc0;
			7784: dout = 12'haa0;
			7785: dout = 12'h000;
			7786: dout = 12'h000;
			7787: dout = 12'h000;

			7788: dout = 12'h000;
			7789: dout = 12'h000;
			7790: dout = 12'h000;
			7791: dout = 12'h000;
			7792: dout = 12'h000;
			7793: dout = 12'h000;
			7794: dout = 12'h000;
			7795: dout = 12'h000;
			7796: dout = 12'h352;
			7797: dout = 12'h883;
			7798: dout = 12'hfc0;
			7799: dout = 12'h550;
			7800: dout = 12'h220;
			7801: dout = 12'h000;
			7802: dout = 12'h000;
			7803: dout = 12'h000;

			7804: dout = 12'h000;
			7805: dout = 12'h000;
			7806: dout = 12'h000;
			7807: dout = 12'h000;
			7808: dout = 12'h000;
			7809: dout = 12'h000;
			7810: dout = 12'h000;
			7811: dout = 12'h011;
			7812: dout = 12'h132;
			7813: dout = 12'h452;
			7814: dout = 12'hbb0;
			7815: dout = 12'h220;
			7816: dout = 12'h110;
			7817: dout = 12'h440;
			7818: dout = 12'h000;
			7819: dout = 12'h000;

			7820: dout = 12'h000;
			7821: dout = 12'h000;
			7822: dout = 12'h000;
			7823: dout = 12'h000;
			7824: dout = 12'h000;
			7825: dout = 12'h000;
			7826: dout = 12'h000;
			7827: dout = 12'h354;
			7828: dout = 12'h011;
			7829: dout = 12'h000;
			7830: dout = 12'h000;
			7831: dout = 12'h000;
			7832: dout = 12'h550;
			7833: dout = 12'hff0;
			7834: dout = 12'h110;
			7835: dout = 12'h000;

			7836: dout = 12'h000;
			7837: dout = 12'h000;
			7838: dout = 12'h000;
			7839: dout = 12'h000;
			7840: dout = 12'h000;
			7841: dout = 12'h000;
			7842: dout = 12'h000;
			7843: dout = 12'h354;
			7844: dout = 12'h011;
			7845: dout = 12'h000;
			7846: dout = 12'h000;
			7847: dout = 12'h000;
			7848: dout = 12'h110;
			7849: dout = 12'h340;
			7850: dout = 12'h000;
			7851: dout = 12'h000;

			7852: dout = 12'h000;
			7853: dout = 12'h000;
			7854: dout = 12'h000;
			7855: dout = 12'h000;
			7856: dout = 12'h011;
			7857: dout = 12'h011;
			7858: dout = 12'h011;
			7859: dout = 12'h254;
			7860: dout = 12'h122;
			7861: dout = 12'h011;
			7862: dout = 12'h011;
			7863: dout = 12'h000;
			7864: dout = 12'h000;
			7865: dout = 12'h000;
			7866: dout = 12'h000;
			7867: dout = 12'h000;

			7868: dout = 12'h000;
			7869: dout = 12'h000;
			7870: dout = 12'h000;
			7871: dout = 12'h000;
			7872: dout = 12'h244;
			7873: dout = 12'h244;
			7874: dout = 12'h244;
			7875: dout = 12'h244;
			7876: dout = 12'h244;
			7877: dout = 12'h244;
			7878: dout = 12'h244;
			7879: dout = 12'h001;
			7880: dout = 12'h000;
			7881: dout = 12'h000;
			7882: dout = 12'h000;
			7883: dout = 12'h000;

			7884: dout = 12'h000;
			7885: dout = 12'h000;
			7886: dout = 12'h011;
			7887: dout = 12'h133;
			7888: dout = 12'h244;
			7889: dout = 12'h244;
			7890: dout = 12'h244;
			7891: dout = 12'h244;
			7892: dout = 12'h89a;
			7893: dout = 12'h9aa;
			7894: dout = 12'h244;
			7895: dout = 12'h133;
			7896: dout = 12'h122;
			7897: dout = 12'h000;
			7898: dout = 12'h000;
			7899: dout = 12'h000;

			7900: dout = 12'h000;
			7901: dout = 12'h000;
			7902: dout = 12'h123;
			7903: dout = 12'h244;
			7904: dout = 12'h244;
			7905: dout = 12'h244;
			7906: dout = 12'h244;
			7907: dout = 12'h244;
			7908: dout = 12'habb;
			7909: dout = 12'hbbb;
			7910: dout = 12'h466;
			7911: dout = 12'h245;
			7912: dout = 12'h133;
			7913: dout = 12'h000;
			7914: dout = 12'h000;
			7915: dout = 12'h000;

			7916: dout = 12'h000;
			7917: dout = 12'h244;
			7918: dout = 12'h244;
			7919: dout = 12'h244;
			7920: dout = 12'h244;
			7921: dout = 12'h244;
			7922: dout = 12'h244;
			7923: dout = 12'h244;
			7924: dout = 12'h244;
			7925: dout = 12'h577;
			7926: dout = 12'hfff;
			7927: dout = 12'h567;
			7928: dout = 12'h244;
			7929: dout = 12'h244;
			7930: dout = 12'h000;
			7931: dout = 12'h000;

			7932: dout = 12'h000;
			7933: dout = 12'h234;
			7934: dout = 12'h244;
			7935: dout = 12'h244;
			7936: dout = 12'h244;
			7937: dout = 12'h244;
			7938: dout = 12'h244;
			7939: dout = 12'h244;
			7940: dout = 12'h244;
			7941: dout = 12'h355;
			7942: dout = 12'h788;
			7943: dout = 12'haab;
			7944: dout = 12'h799;
			7945: dout = 12'h244;
			7946: dout = 12'h000;
			7947: dout = 12'h000;

			7948: dout = 12'h000;
			7949: dout = 12'h133;
			7950: dout = 12'h234;
			7951: dout = 12'h244;
			7952: dout = 12'h244;
			7953: dout = 12'h244;
			7954: dout = 12'h244;
			7955: dout = 12'h244;
			7956: dout = 12'h244;
			7957: dout = 12'h244;
			7958: dout = 12'h244;
			7959: dout = 12'hcdd;
			7960: dout = 12'habb;
			7961: dout = 12'h244;
			7962: dout = 12'h000;
			7963: dout = 12'h000;

			7964: dout = 12'h000;
			7965: dout = 12'h133;
			7966: dout = 12'h234;
			7967: dout = 12'h244;
			7968: dout = 12'h244;
			7969: dout = 12'h244;
			7970: dout = 12'h244;
			7971: dout = 12'h244;
			7972: dout = 12'h244;
			7973: dout = 12'h244;
			7974: dout = 12'h244;
			7975: dout = 12'hcdd;
			7976: dout = 12'habb;
			7977: dout = 12'h244;
			7978: dout = 12'h000;
			7979: dout = 12'h000;

			7980: dout = 12'h000;
			7981: dout = 12'h133;
			7982: dout = 12'h234;
			7983: dout = 12'h234;
			7984: dout = 12'h244;
			7985: dout = 12'h244;
			7986: dout = 12'h244;
			7987: dout = 12'h244;
			7988: dout = 12'h244;
			7989: dout = 12'h244;
			7990: dout = 12'h244;
			7991: dout = 12'h688;
			7992: dout = 12'h677;
			7993: dout = 12'h244;
			7994: dout = 12'h000;
			7995: dout = 12'h000;

			7996: dout = 12'h000;
			7997: dout = 12'h133;
			7998: dout = 12'h133;
			7999: dout = 12'h133;
			8000: dout = 12'h244;
			8001: dout = 12'h244;
			8002: dout = 12'h244;
			8003: dout = 12'h244;
			8004: dout = 12'h244;
			8005: dout = 12'h244;
			8006: dout = 12'h244;
			8007: dout = 12'h244;
			8008: dout = 12'h244;
			8009: dout = 12'h244;
			8010: dout = 12'h000;
			8011: dout = 12'h000;

			8012: dout = 12'h000;
			8013: dout = 12'h133;
			8014: dout = 12'h133;
			8015: dout = 12'h133;
			8016: dout = 12'h133;
			8017: dout = 12'h244;
			8018: dout = 12'h244;
			8019: dout = 12'h244;
			8020: dout = 12'h244;
			8021: dout = 12'h244;
			8022: dout = 12'h244;
			8023: dout = 12'h244;
			8024: dout = 12'h244;
			8025: dout = 12'h244;
			8026: dout = 12'h000;
			8027: dout = 12'h000;

			8028: dout = 12'h000;
			8029: dout = 12'h011;
			8030: dout = 12'h122;
			8031: dout = 12'h133;
			8032: dout = 12'h133;
			8033: dout = 12'h234;
			8034: dout = 12'h234;
			8035: dout = 12'h234;
			8036: dout = 12'h244;
			8037: dout = 12'h244;
			8038: dout = 12'h244;
			8039: dout = 12'h244;
			8040: dout = 12'h234;
			8041: dout = 12'h122;
			8042: dout = 12'h000;
			8043: dout = 12'h000;

			8044: dout = 12'h000;
			8045: dout = 12'h000;
			8046: dout = 12'h111;
			8047: dout = 12'h133;
			8048: dout = 12'h133;
			8049: dout = 12'h133;
			8050: dout = 12'h133;
			8051: dout = 12'h133;
			8052: dout = 12'h244;
			8053: dout = 12'h244;
			8054: dout = 12'h244;
			8055: dout = 12'h244;
			8056: dout = 12'h123;
			8057: dout = 12'h000;
			8058: dout = 12'h000;
			8059: dout = 12'h000;

			8060: dout = 12'h000;
			8061: dout = 12'h000;
			8062: dout = 12'h000;
			8063: dout = 12'h000;
			8064: dout = 12'h133;
			8065: dout = 12'h133;
			8066: dout = 12'h133;
			8067: dout = 12'h133;
			8068: dout = 12'h133;
			8069: dout = 12'h133;
			8070: dout = 12'h133;
			8071: dout = 12'h000;
			8072: dout = 12'h000;
			8073: dout = 12'h000;
			8074: dout = 12'h000;
			8075: dout = 12'h000;

			8076: dout = 12'h000;
			8077: dout = 12'h000;
			8078: dout = 12'h000;
			8079: dout = 12'h000;
			8080: dout = 12'h112;
			8081: dout = 12'h112;
			8082: dout = 12'h112;
			8083: dout = 12'h112;
			8084: dout = 12'h112;
			8085: dout = 12'h112;
			8086: dout = 12'h112;
			8087: dout = 12'h000;
			8088: dout = 12'h000;
			8089: dout = 12'h000;
			8090: dout = 12'h000;
			8091: dout = 12'h000;

			8092: dout = 12'h000;
			8093: dout = 12'h000;
			8094: dout = 12'h000;
			8095: dout = 12'h000;
			8096: dout = 12'h000;
			8097: dout = 12'h000;
			8098: dout = 12'h000;
			8099: dout = 12'h000;
			8100: dout = 12'h000;
			8101: dout = 12'h000;
			8102: dout = 12'h000;
			8103: dout = 12'h000;
			8104: dout = 12'h000;
			8105: dout = 12'h000;
			8106: dout = 12'h000;
			8107: dout = 12'h000;

			8108: dout = 12'h000;
			8109: dout = 12'h000;
			8110: dout = 12'h000;
			8111: dout = 12'h000;
			8112: dout = 12'h000;
			8113: dout = 12'h000;
			8114: dout = 12'h000;
			8115: dout = 12'h000;
			8116: dout = 12'h000;
			8117: dout = 12'h000;
			8118: dout = 12'h000;
			8119: dout = 12'h000;
			8120: dout = 12'h000;
			8121: dout = 12'h000;
			8122: dout = 12'h000;
			8123: dout = 12'h000;

			8124: dout = 12'h000;
			8125: dout = 12'h000;
			8126: dout = 12'h000;
			8127: dout = 12'h000;
			8128: dout = 12'h000;
			8129: dout = 12'h000;
			8130: dout = 12'h000;
			8131: dout = 12'h330;
			8132: dout = 12'h000;
			8133: dout = 12'h000;
			8134: dout = 12'h000;
			8135: dout = 12'h000;
			8136: dout = 12'h000;
			8137: dout = 12'h000;
			8138: dout = 12'h000;
			8139: dout = 12'h000;

			8140: dout = 12'h000;
			8141: dout = 12'h000;
			8142: dout = 12'h000;
			8143: dout = 12'h000;
			8144: dout = 12'h000;
			8145: dout = 12'h000;
			8146: dout = 12'h220;
			8147: dout = 12'hfe0;
			8148: dout = 12'h330;
			8149: dout = 12'h540;
			8150: dout = 12'h500;
			8151: dout = 12'h100;
			8152: dout = 12'h000;
			8153: dout = 12'h000;
			8154: dout = 12'h000;
			8155: dout = 12'h000;

			8156: dout = 12'h000;
			8157: dout = 12'h000;
			8158: dout = 12'h000;
			8159: dout = 12'h000;
			8160: dout = 12'h000;
			8161: dout = 12'h000;
			8162: dout = 12'h000;
			8163: dout = 12'h000;
			8164: dout = 12'hab0;
			8165: dout = 12'hfc0;
			8166: dout = 12'hf00;
			8167: dout = 12'h300;
			8168: dout = 12'h000;
			8169: dout = 12'h000;
			8170: dout = 12'h000;
			8171: dout = 12'h000;

			8172: dout = 12'h000;
			8173: dout = 12'h000;
			8174: dout = 12'h000;
			8175: dout = 12'h000;
			8176: dout = 12'h000;
			8177: dout = 12'h000;
			8178: dout = 12'h000;
			8179: dout = 12'h000;
			8180: dout = 12'h352;
			8181: dout = 12'h883;
			8182: dout = 12'hfc0;
			8183: dout = 12'h320;
			8184: dout = 12'h000;
			8185: dout = 12'h000;
			8186: dout = 12'h000;
			8187: dout = 12'h000;

			8188: dout = 12'h000;
			8189: dout = 12'h000;
			8190: dout = 12'h000;
			8191: dout = 12'h000;
			8192: dout = 12'h000;
			8193: dout = 12'h000;
			8194: dout = 12'h000;
			8195: dout = 12'h011;
			8196: dout = 12'h132;
			8197: dout = 12'h452;
			8198: dout = 12'hbb0;
			8199: dout = 12'h990;
			8200: dout = 12'h980;
			8201: dout = 12'h000;
			8202: dout = 12'h000;
			8203: dout = 12'h000;

			8204: dout = 12'h000;
			8205: dout = 12'h000;
			8206: dout = 12'h000;
			8207: dout = 12'h000;
			8208: dout = 12'h000;
			8209: dout = 12'h000;
			8210: dout = 12'h000;
			8211: dout = 12'h354;
			8212: dout = 12'h011;
			8213: dout = 12'h000;
			8214: dout = 12'h000;
			8215: dout = 12'h220;
			8216: dout = 12'h330;
			8217: dout = 12'h000;
			8218: dout = 12'h000;
			8219: dout = 12'h000;

			8220: dout = 12'h000;
			8221: dout = 12'h000;
			8222: dout = 12'h000;
			8223: dout = 12'h000;
			8224: dout = 12'h000;
			8225: dout = 12'h000;
			8226: dout = 12'h000;
			8227: dout = 12'h354;
			8228: dout = 12'h011;
			8229: dout = 12'h000;
			8230: dout = 12'h000;
			8231: dout = 12'h000;
			8232: dout = 12'h000;
			8233: dout = 12'h000;
			8234: dout = 12'h000;
			8235: dout = 12'h000;

			8236: dout = 12'h000;
			8237: dout = 12'h000;
			8238: dout = 12'h000;
			8239: dout = 12'h000;
			8240: dout = 12'h011;
			8241: dout = 12'h011;
			8242: dout = 12'h011;
			8243: dout = 12'h254;
			8244: dout = 12'h122;
			8245: dout = 12'h011;
			8246: dout = 12'h011;
			8247: dout = 12'h000;
			8248: dout = 12'h000;
			8249: dout = 12'h000;
			8250: dout = 12'h000;
			8251: dout = 12'h000;

			8252: dout = 12'h000;
			8253: dout = 12'h000;
			8254: dout = 12'h000;
			8255: dout = 12'h000;
			8256: dout = 12'h244;
			8257: dout = 12'h244;
			8258: dout = 12'h244;
			8259: dout = 12'h244;
			8260: dout = 12'h244;
			8261: dout = 12'h244;
			8262: dout = 12'h244;
			8263: dout = 12'h001;
			8264: dout = 12'h000;
			8265: dout = 12'h000;
			8266: dout = 12'h000;
			8267: dout = 12'h000;

			8268: dout = 12'h000;
			8269: dout = 12'h000;
			8270: dout = 12'h011;
			8271: dout = 12'h133;
			8272: dout = 12'h244;
			8273: dout = 12'h244;
			8274: dout = 12'h244;
			8275: dout = 12'h244;
			8276: dout = 12'h89a;
			8277: dout = 12'h9aa;
			8278: dout = 12'h244;
			8279: dout = 12'h133;
			8280: dout = 12'h122;
			8281: dout = 12'h000;
			8282: dout = 12'h000;
			8283: dout = 12'h000;

			8284: dout = 12'h000;
			8285: dout = 12'h000;
			8286: dout = 12'h123;
			8287: dout = 12'h244;
			8288: dout = 12'h244;
			8289: dout = 12'h244;
			8290: dout = 12'h244;
			8291: dout = 12'h244;
			8292: dout = 12'habb;
			8293: dout = 12'hbbb;
			8294: dout = 12'h466;
			8295: dout = 12'h245;
			8296: dout = 12'h133;
			8297: dout = 12'h000;
			8298: dout = 12'h000;
			8299: dout = 12'h000;

			8300: dout = 12'h000;
			8301: dout = 12'h244;
			8302: dout = 12'h244;
			8303: dout = 12'h244;
			8304: dout = 12'h244;
			8305: dout = 12'h244;
			8306: dout = 12'h244;
			8307: dout = 12'h244;
			8308: dout = 12'h244;
			8309: dout = 12'h577;
			8310: dout = 12'hfff;
			8311: dout = 12'h567;
			8312: dout = 12'h244;
			8313: dout = 12'h244;
			8314: dout = 12'h000;
			8315: dout = 12'h000;

			8316: dout = 12'h000;
			8317: dout = 12'h234;
			8318: dout = 12'h244;
			8319: dout = 12'h244;
			8320: dout = 12'h244;
			8321: dout = 12'h244;
			8322: dout = 12'h244;
			8323: dout = 12'h244;
			8324: dout = 12'h244;
			8325: dout = 12'h355;
			8326: dout = 12'h788;
			8327: dout = 12'haab;
			8328: dout = 12'h799;
			8329: dout = 12'h244;
			8330: dout = 12'h000;
			8331: dout = 12'h000;

			8332: dout = 12'h000;
			8333: dout = 12'h133;
			8334: dout = 12'h234;
			8335: dout = 12'h244;
			8336: dout = 12'h244;
			8337: dout = 12'h244;
			8338: dout = 12'h244;
			8339: dout = 12'h244;
			8340: dout = 12'h244;
			8341: dout = 12'h244;
			8342: dout = 12'h244;
			8343: dout = 12'hcdd;
			8344: dout = 12'habb;
			8345: dout = 12'h244;
			8346: dout = 12'h000;
			8347: dout = 12'h000;

			8348: dout = 12'h000;
			8349: dout = 12'h133;
			8350: dout = 12'h234;
			8351: dout = 12'h244;
			8352: dout = 12'h244;
			8353: dout = 12'h244;
			8354: dout = 12'h244;
			8355: dout = 12'h244;
			8356: dout = 12'h244;
			8357: dout = 12'h244;
			8358: dout = 12'h244;
			8359: dout = 12'hcdd;
			8360: dout = 12'habb;
			8361: dout = 12'h244;
			8362: dout = 12'h000;
			8363: dout = 12'h000;

			8364: dout = 12'h000;
			8365: dout = 12'h133;
			8366: dout = 12'h234;
			8367: dout = 12'h234;
			8368: dout = 12'h244;
			8369: dout = 12'h244;
			8370: dout = 12'h244;
			8371: dout = 12'h244;
			8372: dout = 12'h244;
			8373: dout = 12'h244;
			8374: dout = 12'h244;
			8375: dout = 12'h688;
			8376: dout = 12'h677;
			8377: dout = 12'h244;
			8378: dout = 12'h000;
			8379: dout = 12'h000;

			8380: dout = 12'h000;
			8381: dout = 12'h133;
			8382: dout = 12'h133;
			8383: dout = 12'h133;
			8384: dout = 12'h244;
			8385: dout = 12'h244;
			8386: dout = 12'h244;
			8387: dout = 12'h244;
			8388: dout = 12'h244;
			8389: dout = 12'h244;
			8390: dout = 12'h244;
			8391: dout = 12'h244;
			8392: dout = 12'h244;
			8393: dout = 12'h244;
			8394: dout = 12'h000;
			8395: dout = 12'h000;

			8396: dout = 12'h000;
			8397: dout = 12'h133;
			8398: dout = 12'h133;
			8399: dout = 12'h133;
			8400: dout = 12'h133;
			8401: dout = 12'h244;
			8402: dout = 12'h244;
			8403: dout = 12'h244;
			8404: dout = 12'h244;
			8405: dout = 12'h244;
			8406: dout = 12'h244;
			8407: dout = 12'h244;
			8408: dout = 12'h244;
			8409: dout = 12'h244;
			8410: dout = 12'h000;
			8411: dout = 12'h000;

			8412: dout = 12'h000;
			8413: dout = 12'h011;
			8414: dout = 12'h122;
			8415: dout = 12'h133;
			8416: dout = 12'h133;
			8417: dout = 12'h234;
			8418: dout = 12'h234;
			8419: dout = 12'h234;
			8420: dout = 12'h244;
			8421: dout = 12'h244;
			8422: dout = 12'h244;
			8423: dout = 12'h244;
			8424: dout = 12'h234;
			8425: dout = 12'h122;
			8426: dout = 12'h000;
			8427: dout = 12'h000;

			8428: dout = 12'h000;
			8429: dout = 12'h000;
			8430: dout = 12'h111;
			8431: dout = 12'h133;
			8432: dout = 12'h133;
			8433: dout = 12'h133;
			8434: dout = 12'h133;
			8435: dout = 12'h133;
			8436: dout = 12'h244;
			8437: dout = 12'h244;
			8438: dout = 12'h244;
			8439: dout = 12'h244;
			8440: dout = 12'h123;
			8441: dout = 12'h000;
			8442: dout = 12'h000;
			8443: dout = 12'h000;

			8444: dout = 12'h000;
			8445: dout = 12'h000;
			8446: dout = 12'h000;
			8447: dout = 12'h000;
			8448: dout = 12'h133;
			8449: dout = 12'h133;
			8450: dout = 12'h133;
			8451: dout = 12'h133;
			8452: dout = 12'h133;
			8453: dout = 12'h133;
			8454: dout = 12'h133;
			8455: dout = 12'h000;
			8456: dout = 12'h000;
			8457: dout = 12'h000;
			8458: dout = 12'h000;
			8459: dout = 12'h000;

			8460: dout = 12'h000;
			8461: dout = 12'h000;
			8462: dout = 12'h000;
			8463: dout = 12'h000;
			8464: dout = 12'h112;
			8465: dout = 12'h112;
			8466: dout = 12'h112;
			8467: dout = 12'h112;
			8468: dout = 12'h112;
			8469: dout = 12'h112;
			8470: dout = 12'h112;
			8471: dout = 12'h000;
			8472: dout = 12'h000;
			8473: dout = 12'h000;
			8474: dout = 12'h000;
			8475: dout = 12'h000;

			8476: dout = 12'h643;
			8477: dout = 12'h521;
			8478: dout = 12'h521;
			8479: dout = 12'h521;
			8480: dout = 12'h521;
			8481: dout = 12'h521;
			8482: dout = 12'h744;
			8483: dout = 12'he87;
			8484: dout = 12'he86;
			8485: dout = 12'he86;
			8486: dout = 12'ha75;
			8487: dout = 12'h643;
			8488: dout = 12'h521;
			8489: dout = 12'h521;
			8490: dout = 12'h521;
			8491: dout = 12'h521;
			8492: dout = 12'h521;
			8493: dout = 12'h644;
			8494: dout = 12'he97;
			8495: dout = 12'he86;
			8496: dout = 12'he86;
			8497: dout = 12'ha75;
			8498: dout = 12'h643;
			8499: dout = 12'h521;
			8500: dout = 12'h521;
			8501: dout = 12'h521;
			8502: dout = 12'h521;
			8503: dout = 12'h521;
			8504: dout = 12'h644;
			8505: dout = 12'he97;
			8506: dout = 12'he86;
			8507: dout = 12'he86;
			8508: dout = 12'ha75;
			8509: dout = 12'h643;
			8510: dout = 12'h521;
			8511: dout = 12'h521;
			8512: dout = 12'h521;
			8513: dout = 12'h521;
			8514: dout = 12'h521;
			8515: dout = 12'h754;
			8516: dout = 12'he97;
			8517: dout = 12'he86;
			8518: dout = 12'he86;
			8519: dout = 12'ha75;
			8520: dout = 12'h643;
			8521: dout = 12'h521;
			8522: dout = 12'h521;
			8523: dout = 12'h521;
			8524: dout = 12'h521;
			8525: dout = 12'h521;
			8526: dout = 12'h754;
			8527: dout = 12'he97;
			8528: dout = 12'he86;
			8529: dout = 12'he86;
			8530: dout = 12'ha65;

			8531: dout = 12'he87;
			8532: dout = 12'hc42;
			8533: dout = 12'hc42;
			8534: dout = 12'hc42;
			8535: dout = 12'hc42;
			8536: dout = 12'ha42;
			8537: dout = 12'h654;
			8538: dout = 12'hd64;
			8539: dout = 12'hc42;
			8540: dout = 12'hc42;
			8541: dout = 12'h411;
			8542: dout = 12'he97;
			8543: dout = 12'hc42;
			8544: dout = 12'hc42;
			8545: dout = 12'hc42;
			8546: dout = 12'hc42;
			8547: dout = 12'ha42;
			8548: dout = 12'h654;
			8549: dout = 12'hd64;
			8550: dout = 12'hc42;
			8551: dout = 12'hc42;
			8552: dout = 12'h411;
			8553: dout = 12'he97;
			8554: dout = 12'hc42;
			8555: dout = 12'hc42;
			8556: dout = 12'hc42;
			8557: dout = 12'hc42;
			8558: dout = 12'ha42;
			8559: dout = 12'h654;
			8560: dout = 12'hd64;
			8561: dout = 12'hc42;
			8562: dout = 12'hc42;
			8563: dout = 12'h411;
			8564: dout = 12'he97;
			8565: dout = 12'hc42;
			8566: dout = 12'hc42;
			8567: dout = 12'hc42;
			8568: dout = 12'hc42;
			8569: dout = 12'ha42;
			8570: dout = 12'h754;
			8571: dout = 12'hd64;
			8572: dout = 12'hc42;
			8573: dout = 12'hc42;
			8574: dout = 12'h410;
			8575: dout = 12'he97;
			8576: dout = 12'hc42;
			8577: dout = 12'hc42;
			8578: dout = 12'hc42;
			8579: dout = 12'hc42;
			8580: dout = 12'ha42;
			8581: dout = 12'h754;
			8582: dout = 12'hd64;
			8583: dout = 12'hc42;
			8584: dout = 12'hc42;
			8585: dout = 12'h421;

			8586: dout = 12'he87;
			8587: dout = 12'hc42;
			8588: dout = 12'hc42;
			8589: dout = 12'hc42;
			8590: dout = 12'hc42;
			8591: dout = 12'ha42;
			8592: dout = 12'h654;
			8593: dout = 12'hd64;
			8594: dout = 12'hc42;
			8595: dout = 12'hc42;
			8596: dout = 12'h411;
			8597: dout = 12'he97;
			8598: dout = 12'hc42;
			8599: dout = 12'hc42;
			8600: dout = 12'hc42;
			8601: dout = 12'hc42;
			8602: dout = 12'ha42;
			8603: dout = 12'h654;
			8604: dout = 12'hd64;
			8605: dout = 12'hc42;
			8606: dout = 12'hc42;
			8607: dout = 12'h411;
			8608: dout = 12'he97;
			8609: dout = 12'hc42;
			8610: dout = 12'hc42;
			8611: dout = 12'hc42;
			8612: dout = 12'hc42;
			8613: dout = 12'ha42;
			8614: dout = 12'h654;
			8615: dout = 12'hd64;
			8616: dout = 12'hc42;
			8617: dout = 12'hc42;
			8618: dout = 12'h411;
			8619: dout = 12'he97;
			8620: dout = 12'hc42;
			8621: dout = 12'hc42;
			8622: dout = 12'hc42;
			8623: dout = 12'hc42;
			8624: dout = 12'ha42;
			8625: dout = 12'h754;
			8626: dout = 12'hd64;
			8627: dout = 12'hc42;
			8628: dout = 12'hc42;
			8629: dout = 12'h411;
			8630: dout = 12'he97;
			8631: dout = 12'hc42;
			8632: dout = 12'hc42;
			8633: dout = 12'hc42;
			8634: dout = 12'hc42;
			8635: dout = 12'ha42;
			8636: dout = 12'h754;
			8637: dout = 12'hd64;
			8638: dout = 12'hc42;
			8639: dout = 12'hc42;
			8640: dout = 12'h421;

			8641: dout = 12'he87;
			8642: dout = 12'hc42;
			8643: dout = 12'hc42;
			8644: dout = 12'hc42;
			8645: dout = 12'hc42;
			8646: dout = 12'ha42;
			8647: dout = 12'h422;
			8648: dout = 12'hb53;
			8649: dout = 12'hc42;
			8650: dout = 12'hc42;
			8651: dout = 12'h411;
			8652: dout = 12'he97;
			8653: dout = 12'hc42;
			8654: dout = 12'hc42;
			8655: dout = 12'hc42;
			8656: dout = 12'hc42;
			8657: dout = 12'ha42;
			8658: dout = 12'h422;
			8659: dout = 12'hb53;
			8660: dout = 12'hc42;
			8661: dout = 12'hc42;
			8662: dout = 12'h411;
			8663: dout = 12'he97;
			8664: dout = 12'hc42;
			8665: dout = 12'hc42;
			8666: dout = 12'hc42;
			8667: dout = 12'hc42;
			8668: dout = 12'ha42;
			8669: dout = 12'h422;
			8670: dout = 12'hb53;
			8671: dout = 12'hc42;
			8672: dout = 12'hc42;
			8673: dout = 12'h411;
			8674: dout = 12'he97;
			8675: dout = 12'hc42;
			8676: dout = 12'hc42;
			8677: dout = 12'hc42;
			8678: dout = 12'hc42;
			8679: dout = 12'ha42;
			8680: dout = 12'h422;
			8681: dout = 12'hb53;
			8682: dout = 12'hc42;
			8683: dout = 12'hc42;
			8684: dout = 12'h411;
			8685: dout = 12'he97;
			8686: dout = 12'hc42;
			8687: dout = 12'hc42;
			8688: dout = 12'hc42;
			8689: dout = 12'hc42;
			8690: dout = 12'ha42;
			8691: dout = 12'h422;
			8692: dout = 12'hb53;
			8693: dout = 12'hc42;
			8694: dout = 12'hc42;
			8695: dout = 12'h421;

			8696: dout = 12'he87;
			8697: dout = 12'hc42;
			8698: dout = 12'hc42;
			8699: dout = 12'hc42;
			8700: dout = 12'hc42;
			8701: dout = 12'h632;
			8702: dout = 12'h654;
			8703: dout = 12'h311;
			8704: dout = 12'h421;
			8705: dout = 12'h421;
			8706: dout = 12'h210;
			8707: dout = 12'he97;
			8708: dout = 12'hc42;
			8709: dout = 12'hc42;
			8710: dout = 12'hc42;
			8711: dout = 12'hc42;
			8712: dout = 12'h632;
			8713: dout = 12'h654;
			8714: dout = 12'h311;
			8715: dout = 12'h421;
			8716: dout = 12'h421;
			8717: dout = 12'h210;
			8718: dout = 12'he97;
			8719: dout = 12'hc42;
			8720: dout = 12'hc42;
			8721: dout = 12'hc42;
			8722: dout = 12'hc42;
			8723: dout = 12'h632;
			8724: dout = 12'h654;
			8725: dout = 12'h311;
			8726: dout = 12'h421;
			8727: dout = 12'h421;
			8728: dout = 12'h210;
			8729: dout = 12'he97;
			8730: dout = 12'hc42;
			8731: dout = 12'hc42;
			8732: dout = 12'hc42;
			8733: dout = 12'hc42;
			8734: dout = 12'h632;
			8735: dout = 12'h644;
			8736: dout = 12'h311;
			8737: dout = 12'h421;
			8738: dout = 12'h421;
			8739: dout = 12'h200;
			8740: dout = 12'he97;
			8741: dout = 12'hc42;
			8742: dout = 12'hc42;
			8743: dout = 12'hc42;
			8744: dout = 12'hc42;
			8745: dout = 12'h632;
			8746: dout = 12'h654;
			8747: dout = 12'h311;
			8748: dout = 12'h421;
			8749: dout = 12'h421;
			8750: dout = 12'h211;

			8751: dout = 12'he87;
			8752: dout = 12'hc42;
			8753: dout = 12'hc42;
			8754: dout = 12'hc42;
			8755: dout = 12'hc42;
			8756: dout = 12'h422;
			8757: dout = 12'hea8;
			8758: dout = 12'he87;
			8759: dout = 12'he97;
			8760: dout = 12'he87;
			8761: dout = 12'h522;
			8762: dout = 12'he97;
			8763: dout = 12'hc42;
			8764: dout = 12'hc42;
			8765: dout = 12'hc42;
			8766: dout = 12'hc42;
			8767: dout = 12'h422;
			8768: dout = 12'hea8;
			8769: dout = 12'he97;
			8770: dout = 12'he97;
			8771: dout = 12'he87;
			8772: dout = 12'h522;
			8773: dout = 12'he97;
			8774: dout = 12'hc42;
			8775: dout = 12'hc42;
			8776: dout = 12'hc42;
			8777: dout = 12'hc42;
			8778: dout = 12'h422;
			8779: dout = 12'hea8;
			8780: dout = 12'he97;
			8781: dout = 12'he97;
			8782: dout = 12'he87;
			8783: dout = 12'h522;
			8784: dout = 12'he97;
			8785: dout = 12'hc42;
			8786: dout = 12'hc42;
			8787: dout = 12'hc42;
			8788: dout = 12'hc42;
			8789: dout = 12'h422;
			8790: dout = 12'hea8;
			8791: dout = 12'he97;
			8792: dout = 12'he97;
			8793: dout = 12'he87;
			8794: dout = 12'h422;
			8795: dout = 12'he97;
			8796: dout = 12'hc42;
			8797: dout = 12'hc42;
			8798: dout = 12'hc42;
			8799: dout = 12'hc42;
			8800: dout = 12'h422;
			8801: dout = 12'hea8;
			8802: dout = 12'he97;
			8803: dout = 12'he97;
			8804: dout = 12'he87;
			8805: dout = 12'h532;

			8806: dout = 12'h743;
			8807: dout = 12'ha32;
			8808: dout = 12'hd52;
			8809: dout = 12'hd52;
			8810: dout = 12'h931;
			8811: dout = 12'h965;
			8812: dout = 12'hd64;
			8813: dout = 12'hc42;
			8814: dout = 12'hc42;
			8815: dout = 12'hc42;
			8816: dout = 12'h411;
			8817: dout = 12'h743;
			8818: dout = 12'ha31;
			8819: dout = 12'hd52;
			8820: dout = 12'hd52;
			8821: dout = 12'h931;
			8822: dout = 12'h965;
			8823: dout = 12'hd64;
			8824: dout = 12'hc42;
			8825: dout = 12'hc42;
			8826: dout = 12'hc42;
			8827: dout = 12'h411;
			8828: dout = 12'h743;
			8829: dout = 12'h931;
			8830: dout = 12'hd52;
			8831: dout = 12'hc52;
			8832: dout = 12'h831;
			8833: dout = 12'h965;
			8834: dout = 12'hd64;
			8835: dout = 12'hc42;
			8836: dout = 12'hc42;
			8837: dout = 12'hc42;
			8838: dout = 12'h411;
			8839: dout = 12'h743;
			8840: dout = 12'h931;
			8841: dout = 12'hd52;
			8842: dout = 12'hd52;
			8843: dout = 12'h931;
			8844: dout = 12'h965;
			8845: dout = 12'hd64;
			8846: dout = 12'hc42;
			8847: dout = 12'hc42;
			8848: dout = 12'hc42;
			8849: dout = 12'h411;
			8850: dout = 12'h743;
			8851: dout = 12'h931;
			8852: dout = 12'hd52;
			8853: dout = 12'hd52;
			8854: dout = 12'h931;
			8855: dout = 12'h965;
			8856: dout = 12'hd64;
			8857: dout = 12'hc42;
			8858: dout = 12'hc42;
			8859: dout = 12'hc42;
			8860: dout = 12'h411;

			8861: dout = 12'hc87;
			8862: dout = 12'h854;
			8863: dout = 12'h522;
			8864: dout = 12'h522;
			8865: dout = 12'h865;
			8866: dout = 12'hc53;
			8867: dout = 12'hc42;
			8868: dout = 12'hc42;
			8869: dout = 12'hc42;
			8870: dout = 12'hc42;
			8871: dout = 12'h411;
			8872: dout = 12'hd97;
			8873: dout = 12'h854;
			8874: dout = 12'h522;
			8875: dout = 12'h522;
			8876: dout = 12'h865;
			8877: dout = 12'hc53;
			8878: dout = 12'hc42;
			8879: dout = 12'hc42;
			8880: dout = 12'hc42;
			8881: dout = 12'hc42;
			8882: dout = 12'h411;
			8883: dout = 12'hd97;
			8884: dout = 12'h854;
			8885: dout = 12'h522;
			8886: dout = 12'h522;
			8887: dout = 12'h865;
			8888: dout = 12'hc53;
			8889: dout = 12'hc42;
			8890: dout = 12'hc42;
			8891: dout = 12'hc42;
			8892: dout = 12'hc42;
			8893: dout = 12'h411;
			8894: dout = 12'hd97;
			8895: dout = 12'h854;
			8896: dout = 12'h522;
			8897: dout = 12'h522;
			8898: dout = 12'h865;
			8899: dout = 12'hc53;
			8900: dout = 12'hc42;
			8901: dout = 12'hc42;
			8902: dout = 12'hc42;
			8903: dout = 12'hc42;
			8904: dout = 12'h411;
			8905: dout = 12'hd97;
			8906: dout = 12'h854;
			8907: dout = 12'h522;
			8908: dout = 12'h522;
			8909: dout = 12'h865;
			8910: dout = 12'hc53;
			8911: dout = 12'hc42;
			8912: dout = 12'hc42;
			8913: dout = 12'hc42;
			8914: dout = 12'hc42;
			8915: dout = 12'h421;

			8916: dout = 12'hc52;
			8917: dout = 12'hd64;
			8918: dout = 12'hd76;
			8919: dout = 12'hd87;
			8920: dout = 12'h744;
			8921: dout = 12'hb42;
			8922: dout = 12'hc42;
			8923: dout = 12'hc42;
			8924: dout = 12'hc42;
			8925: dout = 12'hc42;
			8926: dout = 12'h411;
			8927: dout = 12'hd52;
			8928: dout = 12'hd64;
			8929: dout = 12'hd76;
			8930: dout = 12'hd87;
			8931: dout = 12'h744;
			8932: dout = 12'hb42;
			8933: dout = 12'hc42;
			8934: dout = 12'hc42;
			8935: dout = 12'hc42;
			8936: dout = 12'hc42;
			8937: dout = 12'h411;
			8938: dout = 12'hd53;
			8939: dout = 12'hd64;
			8940: dout = 12'hd76;
			8941: dout = 12'hd87;
			8942: dout = 12'h744;
			8943: dout = 12'hb42;
			8944: dout = 12'hc42;
			8945: dout = 12'hc42;
			8946: dout = 12'hc42;
			8947: dout = 12'hc42;
			8948: dout = 12'h411;
			8949: dout = 12'hd52;
			8950: dout = 12'hd64;
			8951: dout = 12'hd76;
			8952: dout = 12'hd87;
			8953: dout = 12'h744;
			8954: dout = 12'hb42;
			8955: dout = 12'hc42;
			8956: dout = 12'hc42;
			8957: dout = 12'hc42;
			8958: dout = 12'hc42;
			8959: dout = 12'h411;
			8960: dout = 12'hd53;
			8961: dout = 12'hd64;
			8962: dout = 12'hd76;
			8963: dout = 12'hd87;
			8964: dout = 12'h744;
			8965: dout = 12'hb42;
			8966: dout = 12'hc42;
			8967: dout = 12'hc42;
			8968: dout = 12'hc42;
			8969: dout = 12'hc42;
			8970: dout = 12'h411;

			8971: dout = 12'hc42;
			8972: dout = 12'hc42;
			8973: dout = 12'hc42;
			8974: dout = 12'hc53;
			8975: dout = 12'hb76;
			8976: dout = 12'h621;
			8977: dout = 12'hc42;
			8978: dout = 12'hc42;
			8979: dout = 12'hc42;
			8980: dout = 12'hc42;
			8981: dout = 12'h411;
			8982: dout = 12'hd52;
			8983: dout = 12'hc42;
			8984: dout = 12'hc42;
			8985: dout = 12'hc53;
			8986: dout = 12'hb76;
			8987: dout = 12'h731;
			8988: dout = 12'hc42;
			8989: dout = 12'hc42;
			8990: dout = 12'hc42;
			8991: dout = 12'hc42;
			8992: dout = 12'h411;
			8993: dout = 12'hd52;
			8994: dout = 12'hc42;
			8995: dout = 12'hc42;
			8996: dout = 12'hc53;
			8997: dout = 12'hb76;
			8998: dout = 12'h731;
			8999: dout = 12'hc42;
			9000: dout = 12'hc42;
			9001: dout = 12'hc42;
			9002: dout = 12'hc42;
			9003: dout = 12'h411;
			9004: dout = 12'hd52;
			9005: dout = 12'hc42;
			9006: dout = 12'hc42;
			9007: dout = 12'hc53;
			9008: dout = 12'hb76;
			9009: dout = 12'h631;
			9010: dout = 12'hc42;
			9011: dout = 12'hc42;
			9012: dout = 12'hc42;
			9013: dout = 12'hc42;
			9014: dout = 12'h411;
			9015: dout = 12'hd52;
			9016: dout = 12'hc42;
			9017: dout = 12'hc42;
			9018: dout = 12'hc53;
			9019: dout = 12'hb76;
			9020: dout = 12'h731;
			9021: dout = 12'hc42;
			9022: dout = 12'hc42;
			9023: dout = 12'hc42;
			9024: dout = 12'hc42;
			9025: dout = 12'h411;

			9026: dout = 12'ha42;
			9027: dout = 12'ha42;
			9028: dout = 12'ha42;
			9029: dout = 12'ha42;
			9030: dout = 12'hb75;
			9031: dout = 12'h211;
			9032: dout = 12'h311;
			9033: dout = 12'h522;
			9034: dout = 12'h522;
			9035: dout = 12'h522;
			9036: dout = 12'h422;
			9037: dout = 12'hb42;
			9038: dout = 12'ha42;
			9039: dout = 12'ha42;
			9040: dout = 12'ha42;
			9041: dout = 12'hb75;
			9042: dout = 12'h211;
			9043: dout = 12'h311;
			9044: dout = 12'h522;
			9045: dout = 12'h522;
			9046: dout = 12'h522;
			9047: dout = 12'h422;
			9048: dout = 12'hb42;
			9049: dout = 12'ha42;
			9050: dout = 12'ha42;
			9051: dout = 12'ha42;
			9052: dout = 12'hb75;
			9053: dout = 12'h211;
			9054: dout = 12'h311;
			9055: dout = 12'h522;
			9056: dout = 12'h522;
			9057: dout = 12'h522;
			9058: dout = 12'h422;
			9059: dout = 12'hb42;
			9060: dout = 12'ha42;
			9061: dout = 12'ha42;
			9062: dout = 12'ha42;
			9063: dout = 12'hb75;
			9064: dout = 12'h211;
			9065: dout = 12'h311;
			9066: dout = 12'h522;
			9067: dout = 12'h522;
			9068: dout = 12'h522;
			9069: dout = 12'h422;
			9070: dout = 12'hb42;
			9071: dout = 12'ha42;
			9072: dout = 12'ha42;
			9073: dout = 12'ha42;
			9074: dout = 12'hb75;
			9075: dout = 12'h311;
			9076: dout = 12'h311;
			9077: dout = 12'h522;
			9078: dout = 12'h522;
			9079: dout = 12'h522;
			9080: dout = 12'h422;

			9081: dout = 12'h643;
			9082: dout = 12'h521;
			9083: dout = 12'h521;
			9084: dout = 12'h521;
			9085: dout = 12'h521;
			9086: dout = 12'h521;
			9087: dout = 12'h754;
			9088: dout = 12'he97;
			9089: dout = 12'he86;
			9090: dout = 12'he86;
			9091: dout = 12'ha76;
			9092: dout = 12'h643;
			9093: dout = 12'h521;
			9094: dout = 12'h521;
			9095: dout = 12'h521;
			9096: dout = 12'h521;
			9097: dout = 12'h521;
			9098: dout = 12'h654;
			9099: dout = 12'he97;
			9100: dout = 12'he86;
			9101: dout = 12'he86;
			9102: dout = 12'ha76;
			9103: dout = 12'h643;
			9104: dout = 12'h521;
			9105: dout = 12'h521;
			9106: dout = 12'h521;
			9107: dout = 12'h521;
			9108: dout = 12'h521;
			9109: dout = 12'h654;
			9110: dout = 12'he97;
			9111: dout = 12'he86;
			9112: dout = 12'he86;
			9113: dout = 12'ha76;
			9114: dout = 12'h643;
			9115: dout = 12'h521;
			9116: dout = 12'h521;
			9117: dout = 12'h521;
			9118: dout = 12'h521;
			9119: dout = 12'h521;
			9120: dout = 12'h754;
			9121: dout = 12'he97;
			9122: dout = 12'he86;
			9123: dout = 12'he86;
			9124: dout = 12'ha76;
			9125: dout = 12'h643;
			9126: dout = 12'h521;
			9127: dout = 12'h521;
			9128: dout = 12'h521;
			9129: dout = 12'h521;
			9130: dout = 12'h521;
			9131: dout = 12'h754;
			9132: dout = 12'he97;
			9133: dout = 12'he86;
			9134: dout = 12'he86;
			9135: dout = 12'ha76;

			9136: dout = 12'he87;
			9137: dout = 12'hc42;
			9138: dout = 12'hc42;
			9139: dout = 12'hc42;
			9140: dout = 12'hc42;
			9141: dout = 12'ha42;
			9142: dout = 12'h654;
			9143: dout = 12'hd64;
			9144: dout = 12'hc42;
			9145: dout = 12'hc42;
			9146: dout = 12'h411;
			9147: dout = 12'he97;
			9148: dout = 12'hc42;
			9149: dout = 12'hc42;
			9150: dout = 12'hc42;
			9151: dout = 12'hc42;
			9152: dout = 12'ha42;
			9153: dout = 12'h654;
			9154: dout = 12'hd64;
			9155: dout = 12'hc42;
			9156: dout = 12'hc42;
			9157: dout = 12'h411;
			9158: dout = 12'he97;
			9159: dout = 12'hc42;
			9160: dout = 12'hc42;
			9161: dout = 12'hc42;
			9162: dout = 12'hc42;
			9163: dout = 12'ha42;
			9164: dout = 12'h654;
			9165: dout = 12'hd64;
			9166: dout = 12'hc42;
			9167: dout = 12'hc42;
			9168: dout = 12'h411;
			9169: dout = 12'he97;
			9170: dout = 12'hc42;
			9171: dout = 12'hc42;
			9172: dout = 12'hc42;
			9173: dout = 12'hc42;
			9174: dout = 12'ha42;
			9175: dout = 12'h754;
			9176: dout = 12'hd64;
			9177: dout = 12'hc42;
			9178: dout = 12'hc42;
			9179: dout = 12'h410;
			9180: dout = 12'he97;
			9181: dout = 12'hc42;
			9182: dout = 12'hc42;
			9183: dout = 12'hc42;
			9184: dout = 12'hc42;
			9185: dout = 12'ha42;
			9186: dout = 12'h754;
			9187: dout = 12'hd64;
			9188: dout = 12'hc42;
			9189: dout = 12'hc42;
			9190: dout = 12'h421;

			9191: dout = 12'he87;
			9192: dout = 12'hc42;
			9193: dout = 12'hc42;
			9194: dout = 12'hc42;
			9195: dout = 12'hc42;
			9196: dout = 12'ha42;
			9197: dout = 12'h654;
			9198: dout = 12'hd64;
			9199: dout = 12'hc42;
			9200: dout = 12'hc42;
			9201: dout = 12'h411;
			9202: dout = 12'he97;
			9203: dout = 12'hc42;
			9204: dout = 12'hc42;
			9205: dout = 12'hc42;
			9206: dout = 12'hc42;
			9207: dout = 12'ha42;
			9208: dout = 12'h654;
			9209: dout = 12'hd64;
			9210: dout = 12'hc42;
			9211: dout = 12'hc42;
			9212: dout = 12'h411;
			9213: dout = 12'he97;
			9214: dout = 12'hc42;
			9215: dout = 12'hc42;
			9216: dout = 12'hc42;
			9217: dout = 12'hc42;
			9218: dout = 12'ha42;
			9219: dout = 12'h654;
			9220: dout = 12'hd64;
			9221: dout = 12'hc42;
			9222: dout = 12'hc42;
			9223: dout = 12'h411;
			9224: dout = 12'he97;
			9225: dout = 12'hc42;
			9226: dout = 12'hc42;
			9227: dout = 12'hc42;
			9228: dout = 12'hc42;
			9229: dout = 12'ha42;
			9230: dout = 12'h754;
			9231: dout = 12'hd64;
			9232: dout = 12'hc42;
			9233: dout = 12'hc42;
			9234: dout = 12'h411;
			9235: dout = 12'he97;
			9236: dout = 12'hc42;
			9237: dout = 12'hc42;
			9238: dout = 12'hc42;
			9239: dout = 12'hc42;
			9240: dout = 12'ha42;
			9241: dout = 12'h754;
			9242: dout = 12'hd64;
			9243: dout = 12'hc42;
			9244: dout = 12'hc42;
			9245: dout = 12'h421;

			9246: dout = 12'he87;
			9247: dout = 12'hc42;
			9248: dout = 12'hc42;
			9249: dout = 12'hc42;
			9250: dout = 12'hc42;
			9251: dout = 12'ha42;
			9252: dout = 12'h422;
			9253: dout = 12'hb53;
			9254: dout = 12'hc42;
			9255: dout = 12'hc42;
			9256: dout = 12'h411;
			9257: dout = 12'he97;
			9258: dout = 12'hc42;
			9259: dout = 12'hc42;
			9260: dout = 12'hc42;
			9261: dout = 12'hc42;
			9262: dout = 12'ha42;
			9263: dout = 12'h322;
			9264: dout = 12'hb53;
			9265: dout = 12'hc42;
			9266: dout = 12'hc42;
			9267: dout = 12'h411;
			9268: dout = 12'he97;
			9269: dout = 12'hc42;
			9270: dout = 12'hc42;
			9271: dout = 12'hc42;
			9272: dout = 12'hc42;
			9273: dout = 12'ha42;
			9274: dout = 12'h322;
			9275: dout = 12'hb53;
			9276: dout = 12'hc42;
			9277: dout = 12'hc42;
			9278: dout = 12'h411;
			9279: dout = 12'he97;
			9280: dout = 12'hc42;
			9281: dout = 12'hc42;
			9282: dout = 12'hc42;
			9283: dout = 12'hc42;
			9284: dout = 12'ha42;
			9285: dout = 12'h422;
			9286: dout = 12'hb53;
			9287: dout = 12'hc42;
			9288: dout = 12'hc42;
			9289: dout = 12'h411;
			9290: dout = 12'he97;
			9291: dout = 12'hc42;
			9292: dout = 12'hc42;
			9293: dout = 12'hc42;
			9294: dout = 12'hc42;
			9295: dout = 12'ha42;
			9296: dout = 12'h422;
			9297: dout = 12'hb53;
			9298: dout = 12'hc42;
			9299: dout = 12'hc42;
			9300: dout = 12'h421;

			9301: dout = 12'he87;
			9302: dout = 12'hc42;
			9303: dout = 12'hc42;
			9304: dout = 12'hc42;
			9305: dout = 12'hc42;
			9306: dout = 12'h632;
			9307: dout = 12'h654;
			9308: dout = 12'h311;
			9309: dout = 12'h421;
			9310: dout = 12'h421;
			9311: dout = 12'h210;
			9312: dout = 12'he97;
			9313: dout = 12'hc42;
			9314: dout = 12'hc42;
			9315: dout = 12'hc42;
			9316: dout = 12'hc42;
			9317: dout = 12'h632;
			9318: dout = 12'h654;
			9319: dout = 12'h311;
			9320: dout = 12'h421;
			9321: dout = 12'h421;
			9322: dout = 12'h210;
			9323: dout = 12'he97;
			9324: dout = 12'hc42;
			9325: dout = 12'hc42;
			9326: dout = 12'hc42;
			9327: dout = 12'hc42;
			9328: dout = 12'h632;
			9329: dout = 12'h754;
			9330: dout = 12'h311;
			9331: dout = 12'h421;
			9332: dout = 12'h421;
			9333: dout = 12'h210;
			9334: dout = 12'he97;
			9335: dout = 12'hc42;
			9336: dout = 12'hc42;
			9337: dout = 12'hc42;
			9338: dout = 12'hc42;
			9339: dout = 12'h632;
			9340: dout = 12'h654;
			9341: dout = 12'h311;
			9342: dout = 12'h421;
			9343: dout = 12'h421;
			9344: dout = 12'h200;
			9345: dout = 12'he97;
			9346: dout = 12'hc42;
			9347: dout = 12'hc42;
			9348: dout = 12'hc42;
			9349: dout = 12'hc42;
			9350: dout = 12'h632;
			9351: dout = 12'h654;
			9352: dout = 12'h311;
			9353: dout = 12'h421;
			9354: dout = 12'h421;
			9355: dout = 12'h211;

			9356: dout = 12'he87;
			9357: dout = 12'hc42;
			9358: dout = 12'hc42;
			9359: dout = 12'hc42;
			9360: dout = 12'hc42;
			9361: dout = 12'h421;
			9362: dout = 12'hea8;
			9363: dout = 12'he97;
			9364: dout = 12'he97;
			9365: dout = 12'he97;
			9366: dout = 12'h522;
			9367: dout = 12'he97;
			9368: dout = 12'hc42;
			9369: dout = 12'hc42;
			9370: dout = 12'hc42;
			9371: dout = 12'hc42;
			9372: dout = 12'h422;
			9373: dout = 12'hea8;
			9374: dout = 12'he97;
			9375: dout = 12'he97;
			9376: dout = 12'he97;
			9377: dout = 12'h522;
			9378: dout = 12'he97;
			9379: dout = 12'hc42;
			9380: dout = 12'hc42;
			9381: dout = 12'hc42;
			9382: dout = 12'hc42;
			9383: dout = 12'h422;
			9384: dout = 12'hea8;
			9385: dout = 12'he97;
			9386: dout = 12'he97;
			9387: dout = 12'he97;
			9388: dout = 12'h522;
			9389: dout = 12'he97;
			9390: dout = 12'hc42;
			9391: dout = 12'hc42;
			9392: dout = 12'hc42;
			9393: dout = 12'hc42;
			9394: dout = 12'h422;
			9395: dout = 12'hea8;
			9396: dout = 12'he97;
			9397: dout = 12'he97;
			9398: dout = 12'he97;
			9399: dout = 12'h422;
			9400: dout = 12'he97;
			9401: dout = 12'hc42;
			9402: dout = 12'hc42;
			9403: dout = 12'hc42;
			9404: dout = 12'hc42;
			9405: dout = 12'h422;
			9406: dout = 12'hea8;
			9407: dout = 12'he97;
			9408: dout = 12'he97;
			9409: dout = 12'he97;
			9410: dout = 12'h532;

			9411: dout = 12'h643;
			9412: dout = 12'h931;
			9413: dout = 12'hc52;
			9414: dout = 12'hc52;
			9415: dout = 12'h831;
			9416: dout = 12'h965;
			9417: dout = 12'hd64;
			9418: dout = 12'hc42;
			9419: dout = 12'hc42;
			9420: dout = 12'hc42;
			9421: dout = 12'h411;
			9422: dout = 12'h743;
			9423: dout = 12'h931;
			9424: dout = 12'hc52;
			9425: dout = 12'hc52;
			9426: dout = 12'h831;
			9427: dout = 12'h965;
			9428: dout = 12'hd64;
			9429: dout = 12'hc42;
			9430: dout = 12'hc42;
			9431: dout = 12'hc42;
			9432: dout = 12'h411;
			9433: dout = 12'h743;
			9434: dout = 12'h931;
			9435: dout = 12'hc52;
			9436: dout = 12'hc52;
			9437: dout = 12'h831;
			9438: dout = 12'h965;
			9439: dout = 12'hd64;
			9440: dout = 12'hc42;
			9441: dout = 12'hc42;
			9442: dout = 12'hc42;
			9443: dout = 12'h411;
			9444: dout = 12'h743;
			9445: dout = 12'h931;
			9446: dout = 12'hc52;
			9447: dout = 12'hc52;
			9448: dout = 12'h831;
			9449: dout = 12'h965;
			9450: dout = 12'hd64;
			9451: dout = 12'hc42;
			9452: dout = 12'hc42;
			9453: dout = 12'hc42;
			9454: dout = 12'h411;
			9455: dout = 12'h743;
			9456: dout = 12'h931;
			9457: dout = 12'hc52;
			9458: dout = 12'hc52;
			9459: dout = 12'h831;
			9460: dout = 12'h965;
			9461: dout = 12'hd64;
			9462: dout = 12'hc42;
			9463: dout = 12'hc42;
			9464: dout = 12'hc42;
			9465: dout = 12'h411;

			9466: dout = 12'hc87;
			9467: dout = 12'h854;
			9468: dout = 12'h532;
			9469: dout = 12'h532;
			9470: dout = 12'h865;
			9471: dout = 12'hc53;
			9472: dout = 12'hc42;
			9473: dout = 12'hc42;
			9474: dout = 12'hc42;
			9475: dout = 12'hc42;
			9476: dout = 12'h411;
			9477: dout = 12'hd97;
			9478: dout = 12'h854;
			9479: dout = 12'h532;
			9480: dout = 12'h532;
			9481: dout = 12'h865;
			9482: dout = 12'hc53;
			9483: dout = 12'hc42;
			9484: dout = 12'hc42;
			9485: dout = 12'hc42;
			9486: dout = 12'hc42;
			9487: dout = 12'h411;
			9488: dout = 12'hd97;
			9489: dout = 12'h854;
			9490: dout = 12'h532;
			9491: dout = 12'h532;
			9492: dout = 12'h865;
			9493: dout = 12'hc53;
			9494: dout = 12'hc42;
			9495: dout = 12'hc42;
			9496: dout = 12'hc42;
			9497: dout = 12'hc42;
			9498: dout = 12'h411;
			9499: dout = 12'hd97;
			9500: dout = 12'h854;
			9501: dout = 12'h532;
			9502: dout = 12'h532;
			9503: dout = 12'h865;
			9504: dout = 12'hc53;
			9505: dout = 12'hc42;
			9506: dout = 12'hc42;
			9507: dout = 12'hc42;
			9508: dout = 12'hc42;
			9509: dout = 12'h411;
			9510: dout = 12'hd97;
			9511: dout = 12'h854;
			9512: dout = 12'h532;
			9513: dout = 12'h532;
			9514: dout = 12'h865;
			9515: dout = 12'hc53;
			9516: dout = 12'hc42;
			9517: dout = 12'hc42;
			9518: dout = 12'hc42;
			9519: dout = 12'hc42;
			9520: dout = 12'h421;

			9521: dout = 12'hc52;
			9522: dout = 12'hd64;
			9523: dout = 12'hd76;
			9524: dout = 12'hd87;
			9525: dout = 12'h744;
			9526: dout = 12'hb42;
			9527: dout = 12'hc42;
			9528: dout = 12'hc42;
			9529: dout = 12'hc42;
			9530: dout = 12'hc42;
			9531: dout = 12'h411;
			9532: dout = 12'hd52;
			9533: dout = 12'hd64;
			9534: dout = 12'hd76;
			9535: dout = 12'hd87;
			9536: dout = 12'h744;
			9537: dout = 12'hb42;
			9538: dout = 12'hc42;
			9539: dout = 12'hc42;
			9540: dout = 12'hc42;
			9541: dout = 12'hc42;
			9542: dout = 12'h411;
			9543: dout = 12'hd52;
			9544: dout = 12'hd64;
			9545: dout = 12'hd76;
			9546: dout = 12'hd87;
			9547: dout = 12'h744;
			9548: dout = 12'hb42;
			9549: dout = 12'hc42;
			9550: dout = 12'hc42;
			9551: dout = 12'hc42;
			9552: dout = 12'hc42;
			9553: dout = 12'h411;
			9554: dout = 12'hd52;
			9555: dout = 12'hd64;
			9556: dout = 12'hd76;
			9557: dout = 12'hd87;
			9558: dout = 12'h744;
			9559: dout = 12'hb42;
			9560: dout = 12'hc42;
			9561: dout = 12'hc42;
			9562: dout = 12'hc42;
			9563: dout = 12'hc42;
			9564: dout = 12'h411;
			9565: dout = 12'hd52;
			9566: dout = 12'hd64;
			9567: dout = 12'hd76;
			9568: dout = 12'hd87;
			9569: dout = 12'h744;
			9570: dout = 12'hb42;
			9571: dout = 12'hc42;
			9572: dout = 12'hc42;
			9573: dout = 12'hc42;
			9574: dout = 12'hc42;
			9575: dout = 12'h411;

			9576: dout = 12'hc42;
			9577: dout = 12'hc42;
			9578: dout = 12'hc42;
			9579: dout = 12'hc53;
			9580: dout = 12'hb76;
			9581: dout = 12'h621;
			9582: dout = 12'hc42;
			9583: dout = 12'hc42;
			9584: dout = 12'hc42;
			9585: dout = 12'hc42;
			9586: dout = 12'h411;
			9587: dout = 12'hd52;
			9588: dout = 12'hc42;
			9589: dout = 12'hc42;
			9590: dout = 12'hc53;
			9591: dout = 12'hb76;
			9592: dout = 12'h621;
			9593: dout = 12'hc42;
			9594: dout = 12'hc42;
			9595: dout = 12'hc42;
			9596: dout = 12'hc42;
			9597: dout = 12'h411;
			9598: dout = 12'hd52;
			9599: dout = 12'hc42;
			9600: dout = 12'hc42;
			9601: dout = 12'hc53;
			9602: dout = 12'hb76;
			9603: dout = 12'h631;
			9604: dout = 12'hc42;
			9605: dout = 12'hc42;
			9606: dout = 12'hc42;
			9607: dout = 12'hc42;
			9608: dout = 12'h411;
			9609: dout = 12'hd52;
			9610: dout = 12'hc42;
			9611: dout = 12'hc42;
			9612: dout = 12'hc53;
			9613: dout = 12'hb76;
			9614: dout = 12'h631;
			9615: dout = 12'hc42;
			9616: dout = 12'hc42;
			9617: dout = 12'hc42;
			9618: dout = 12'hc42;
			9619: dout = 12'h411;
			9620: dout = 12'hd52;
			9621: dout = 12'hc42;
			9622: dout = 12'hc42;
			9623: dout = 12'hc53;
			9624: dout = 12'hb76;
			9625: dout = 12'h631;
			9626: dout = 12'hc42;
			9627: dout = 12'hc42;
			9628: dout = 12'hc42;
			9629: dout = 12'hc42;
			9630: dout = 12'h411;

			9631: dout = 12'ha42;
			9632: dout = 12'ha42;
			9633: dout = 12'ha42;
			9634: dout = 12'ha42;
			9635: dout = 12'hb75;
			9636: dout = 12'h211;
			9637: dout = 12'h211;
			9638: dout = 12'h211;
			9639: dout = 12'h211;
			9640: dout = 12'h211;
			9641: dout = 12'h100;
			9642: dout = 12'ha42;
			9643: dout = 12'ha42;
			9644: dout = 12'ha42;
			9645: dout = 12'ha42;
			9646: dout = 12'hb75;
			9647: dout = 12'h211;
			9648: dout = 12'h211;
			9649: dout = 12'h211;
			9650: dout = 12'h211;
			9651: dout = 12'h211;
			9652: dout = 12'h101;
			9653: dout = 12'ha42;
			9654: dout = 12'ha42;
			9655: dout = 12'ha42;
			9656: dout = 12'ha42;
			9657: dout = 12'hb75;
			9658: dout = 12'h211;
			9659: dout = 12'h211;
			9660: dout = 12'h211;
			9661: dout = 12'h211;
			9662: dout = 12'h211;
			9663: dout = 12'h101;
			9664: dout = 12'ha42;
			9665: dout = 12'ha42;
			9666: dout = 12'ha42;
			9667: dout = 12'ha42;
			9668: dout = 12'hb75;
			9669: dout = 12'h211;
			9670: dout = 12'h211;
			9671: dout = 12'h211;
			9672: dout = 12'h211;
			9673: dout = 12'h211;
			9674: dout = 12'h101;
			9675: dout = 12'ha42;
			9676: dout = 12'ha42;
			9677: dout = 12'ha42;
			9678: dout = 12'ha42;
			9679: dout = 12'hb75;
			9680: dout = 12'h211;
			9681: dout = 12'h211;
			9682: dout = 12'h211;
			9683: dout = 12'h211;
			9684: dout = 12'h211;
			9685: dout = 12'h211;

			9686: dout = 12'h000;
			9687: dout = 12'h000;
			9688: dout = 12'h000;
			9689: dout = 12'h000;
			9690: dout = 12'h000;
			9691: dout = 12'h114;
			9692: dout = 12'h34c;
			9693: dout = 12'h114;
			9694: dout = 12'h000;
			9695: dout = 12'h113;
			9696: dout = 12'h34c;
			9697: dout = 12'h34c;
			9698: dout = 12'h238;
			9699: dout = 12'h002;
			9700: dout = 12'h000;
			9701: dout = 12'h000;
			9702: dout = 12'h000;
			9703: dout = 12'h000;

			9704: dout = 12'h000;
			9705: dout = 12'h000;
			9706: dout = 12'h000;
			9707: dout = 12'h000;
			9708: dout = 12'h115;
			9709: dout = 12'h34a;
			9710: dout = 12'h35a;
			9711: dout = 12'h000;
			9712: dout = 12'h000;
			9713: dout = 12'h258;
			9714: dout = 12'h34a;
			9715: dout = 12'h226;
			9716: dout = 12'h001;
			9717: dout = 12'h237;
			9718: dout = 12'h114;
			9719: dout = 12'h000;
			9720: dout = 12'h000;
			9721: dout = 12'h000;

			9722: dout = 12'h000;
			9723: dout = 12'h000;
			9724: dout = 12'h001;
			9725: dout = 12'h115;
			9726: dout = 12'h34b;
			9727: dout = 12'h46e;
			9728: dout = 12'h36a;
			9729: dout = 12'h000;
			9730: dout = 12'h000;
			9731: dout = 12'h36b;
			9732: dout = 12'h011;
			9733: dout = 12'h458;
			9734: dout = 12'h36b;
			9735: dout = 12'h46e;
			9736: dout = 12'h34a;
			9737: dout = 12'h113;
			9738: dout = 12'h001;
			9739: dout = 12'h000;

			9740: dout = 12'h000;
			9741: dout = 12'h000;
			9742: dout = 12'h113;
			9743: dout = 12'h33a;
			9744: dout = 12'h46c;
			9745: dout = 12'h48e;
			9746: dout = 12'h36a;
			9747: dout = 12'h000;
			9748: dout = 12'h000;
			9749: dout = 12'h000;
			9750: dout = 12'h000;
			9751: dout = 12'h79b;
			9752: dout = 12'h36a;
			9753: dout = 12'h135;
			9754: dout = 12'h012;
			9755: dout = 12'h229;
			9756: dout = 12'h002;
			9757: dout = 12'h000;

			9758: dout = 12'h001;
			9759: dout = 12'h126;
			9760: dout = 12'h236;
			9761: dout = 12'h135;
			9762: dout = 12'h123;
			9763: dout = 12'h247;
			9764: dout = 12'h135;
			9765: dout = 12'h000;
			9766: dout = 12'h000;
			9767: dout = 12'h000;
			9768: dout = 12'h000;
			9769: dout = 12'h345;
			9770: dout = 12'h000;
			9771: dout = 12'h123;
			9772: dout = 12'h47c;
			9773: dout = 12'h247;
			9774: dout = 12'h226;
			9775: dout = 12'h115;

			9776: dout = 12'h001;
			9777: dout = 12'h33a;
			9778: dout = 12'h46d;
			9779: dout = 12'h48d;
			9780: dout = 12'h36a;
			9781: dout = 12'h36a;
			9782: dout = 12'h000;
			9783: dout = 12'h000;
			9784: dout = 12'h000;
			9785: dout = 12'h000;
			9786: dout = 12'h000;
			9787: dout = 12'h000;
			9788: dout = 12'h000;
			9789: dout = 12'h247;
			9790: dout = 12'h48e;
			9791: dout = 12'h48e;
			9792: dout = 12'h238;
			9793: dout = 12'h115;

			9794: dout = 12'h001;
			9795: dout = 12'h339;
			9796: dout = 12'h45d;
			9797: dout = 12'h48e;
			9798: dout = 12'h48e;
			9799: dout = 12'h48e;
			9800: dout = 12'h248;
			9801: dout = 12'h000;
			9802: dout = 12'h000;
			9803: dout = 12'h000;
			9804: dout = 12'h000;
			9805: dout = 12'h000;
			9806: dout = 12'h000;
			9807: dout = 12'h000;
			9808: dout = 12'h000;
			9809: dout = 12'h000;
			9810: dout = 12'h000;
			9811: dout = 12'h114;

			9812: dout = 12'h001;
			9813: dout = 12'h339;
			9814: dout = 12'h45d;
			9815: dout = 12'h48e;
			9816: dout = 12'h36a;
			9817: dout = 12'h247;
			9818: dout = 12'h000;
			9819: dout = 12'h000;
			9820: dout = 12'h000;
			9821: dout = 12'h000;
			9822: dout = 12'h000;
			9823: dout = 12'h000;
			9824: dout = 12'h000;
			9825: dout = 12'h000;
			9826: dout = 12'h000;
			9827: dout = 12'h247;
			9828: dout = 12'h226;
			9829: dout = 12'h125;

			9830: dout = 12'h001;
			9831: dout = 12'h339;
			9832: dout = 12'h125;
			9833: dout = 12'h123;
			9834: dout = 12'h011;
			9835: dout = 12'h000;
			9836: dout = 12'h000;
			9837: dout = 12'h000;
			9838: dout = 12'h000;
			9839: dout = 12'h000;
			9840: dout = 12'h000;
			9841: dout = 12'h000;
			9842: dout = 12'h012;
			9843: dout = 12'h36a;
			9844: dout = 12'h36a;
			9845: dout = 12'h48e;
			9846: dout = 12'h45d;
			9847: dout = 12'h227;

			9848: dout = 12'h001;
			9849: dout = 12'h002;
			9850: dout = 12'h34a;
			9851: dout = 12'h48e;
			9852: dout = 12'h247;
			9853: dout = 12'h000;
			9854: dout = 12'h000;
			9855: dout = 12'h000;
			9856: dout = 12'h000;
			9857: dout = 12'h000;
			9858: dout = 12'h000;
			9859: dout = 12'h248;
			9860: dout = 12'h123;
			9861: dout = 12'h123;
			9862: dout = 12'h123;
			9863: dout = 12'h113;
			9864: dout = 12'h45d;
			9865: dout = 12'h227;

			9866: dout = 12'h000;
			9867: dout = 12'h113;
			9868: dout = 12'h35b;
			9869: dout = 12'h48e;
			9870: dout = 12'h247;
			9871: dout = 12'h135;
			9872: dout = 12'h247;
			9873: dout = 12'h123;
			9874: dout = 12'h000;
			9875: dout = 12'h000;
			9876: dout = 12'h000;
			9877: dout = 12'h000;
			9878: dout = 12'h259;
			9879: dout = 12'h48e;
			9880: dout = 12'h48e;
			9881: dout = 12'h001;
			9882: dout = 12'h33a;
			9883: dout = 12'h227;

			9884: dout = 12'h000;
			9885: dout = 12'h227;
			9886: dout = 12'h46e;
			9887: dout = 12'h48e;
			9888: dout = 12'h247;
			9889: dout = 12'h36a;
			9890: dout = 12'h48e;
			9891: dout = 12'h247;
			9892: dout = 12'h000;
			9893: dout = 12'h000;
			9894: dout = 12'h000;
			9895: dout = 12'h000;
			9896: dout = 12'h123;
			9897: dout = 12'h48e;
			9898: dout = 12'h48e;
			9899: dout = 12'h258;
			9900: dout = 12'h001;
			9901: dout = 12'h115;

			9902: dout = 12'h000;
			9903: dout = 12'h000;
			9904: dout = 12'h114;
			9905: dout = 12'h34c;
			9906: dout = 12'h125;
			9907: dout = 12'h36a;
			9908: dout = 12'h48e;
			9909: dout = 12'h247;
			9910: dout = 12'h248;
			9911: dout = 12'h48e;
			9912: dout = 12'h48e;
			9913: dout = 12'h236;
			9914: dout = 12'h012;
			9915: dout = 12'h135;
			9916: dout = 12'h46c;
			9917: dout = 12'h33b;
			9918: dout = 12'h002;
			9919: dout = 12'h000;

			9920: dout = 12'h000;
			9921: dout = 12'h000;
			9922: dout = 12'h002;
			9923: dout = 12'h114;
			9924: dout = 12'h113;
			9925: dout = 12'h36c;
			9926: dout = 12'h48e;
			9927: dout = 12'h36a;
			9928: dout = 12'h011;
			9929: dout = 12'h259;
			9930: dout = 12'h48e;
			9931: dout = 12'h48e;
			9932: dout = 12'h47c;
			9933: dout = 12'h113;
			9934: dout = 12'h226;
			9935: dout = 12'h114;
			9936: dout = 12'h001;
			9937: dout = 12'h000;

			9938: dout = 12'h000;
			9939: dout = 12'h000;
			9940: dout = 12'h000;
			9941: dout = 12'h000;
			9942: dout = 12'h115;
			9943: dout = 12'h34a;
			9944: dout = 12'h47e;
			9945: dout = 12'h48e;
			9946: dout = 12'h123;
			9947: dout = 12'h000;
			9948: dout = 12'h259;
			9949: dout = 12'h47e;
			9950: dout = 12'h46d;
			9951: dout = 12'h125;
			9952: dout = 12'h113;
			9953: dout = 12'h000;
			9954: dout = 12'h000;
			9955: dout = 12'h000;

			9956: dout = 12'h000;
			9957: dout = 12'h000;
			9958: dout = 12'h000;
			9959: dout = 12'h000;
			9960: dout = 12'h000;
			9961: dout = 12'h113;
			9962: dout = 12'h34b;
			9963: dout = 12'h36b;
			9964: dout = 12'h012;
			9965: dout = 12'h000;
			9966: dout = 12'h247;
			9967: dout = 12'h46d;
			9968: dout = 12'h33a;
			9969: dout = 12'h002;
			9970: dout = 12'h000;
			9971: dout = 12'h000;
			9972: dout = 12'h000;
			9973: dout = 12'h000;

			9974: dout = 12'h000;
			9975: dout = 12'h000;
			9976: dout = 12'h000;
			9977: dout = 12'h000;
			9978: dout = 12'h000;
			9979: dout = 12'h000;
			9980: dout = 12'h002;
			9981: dout = 12'h002;
			9982: dout = 12'h000;
			9983: dout = 12'h000;
			9984: dout = 12'h113;
			9985: dout = 12'h227;
			9986: dout = 12'h001;
			9987: dout = 12'h000;
			9988: dout = 12'h000;
			9989: dout = 12'h000;
			9990: dout = 12'h000;
			9991: dout = 12'h000;

			9992: dout = 12'h000;
			9993: dout = 12'h000;
			9994: dout = 12'h000;
			9995: dout = 12'h000;
			9996: dout = 12'h000;
			9997: dout = 12'h000;
			9998: dout = 12'h000;
			9999: dout = 12'h000;
			10000: dout = 12'h000;
			10001: dout = 12'h001;
			10002: dout = 12'h002;
			10003: dout = 12'h001;
			10004: dout = 12'h000;
			10005: dout = 12'h000;
			10006: dout = 12'h000;
			10007: dout = 12'h000;
			10008: dout = 12'h000;
			10009: dout = 12'h000;

			10010: dout = 12'h000;
			10011: dout = 12'h000;
			10012: dout = 12'h000;
			10013: dout = 12'h000;
			10014: dout = 12'h000;
			10015: dout = 12'h000;
			10016: dout = 12'h000;
			10017: dout = 12'h000;
			10018: dout = 12'h000;
			10019: dout = 12'h001;
			10020: dout = 12'h002;
			10021: dout = 12'h000;
			10022: dout = 12'h000;
			10023: dout = 12'h000;
			10024: dout = 12'h000;
			10025: dout = 12'h000;
			10026: dout = 12'h000;
			10027: dout = 12'h000;

			10028: dout = 12'h000;
			10029: dout = 12'h000;
			10030: dout = 12'h000;
			10031: dout = 12'h000;
			10032: dout = 12'h000;
			10033: dout = 12'h000;
			10034: dout = 12'h000;
			10035: dout = 12'h000;
			10036: dout = 12'h000;
			10037: dout = 12'h000;
			10038: dout = 12'h000;
			10039: dout = 12'h000;
			10040: dout = 12'h000;
			10041: dout = 12'h000;
			10042: dout = 12'h000;
			10043: dout = 12'h000;
			10044: dout = 12'h000;
			10045: dout = 12'h000;

			10046: dout = 12'h000;
			10047: dout = 12'h000;
			10048: dout = 12'h000;
			10049: dout = 12'h000;
			10050: dout = 12'h000;
			10051: dout = 12'h000;
			10052: dout = 12'h000;
			10053: dout = 12'h000;
			10054: dout = 12'h000;
			10055: dout = 12'h000;
			10056: dout = 12'h000;
			10057: dout = 12'h000;
			10058: dout = 12'h000;
			10059: dout = 12'h000;
			10060: dout = 12'h000;
			10061: dout = 12'h000;
			10062: dout = 12'h000;
			10063: dout = 12'h000;

			10064: dout = 12'h000;
			10065: dout = 12'h000;
			10066: dout = 12'h000;
			10067: dout = 12'h000;
			10068: dout = 12'h000;
			10069: dout = 12'h000;
			10070: dout = 12'h000;
			10071: dout = 12'h000;
			10072: dout = 12'h000;
			10073: dout = 12'h000;
			10074: dout = 12'h000;
			10075: dout = 12'h000;
			10076: dout = 12'h000;
			10077: dout = 12'h000;
			10078: dout = 12'h000;
			10079: dout = 12'h000;
			10080: dout = 12'h000;
			10081: dout = 12'h000;

			10082: dout = 12'h000;
			10083: dout = 12'h000;
			10084: dout = 12'h000;
			10085: dout = 12'h000;
			10086: dout = 12'h000;
			10087: dout = 12'h000;
			10088: dout = 12'h000;
			10089: dout = 12'h000;
			10090: dout = 12'h000;
			10091: dout = 12'h000;
			10092: dout = 12'h000;
			10093: dout = 12'h000;
			10094: dout = 12'h000;
			10095: dout = 12'h000;
			10096: dout = 12'h000;
			10097: dout = 12'h000;
			10098: dout = 12'h000;
			10099: dout = 12'h000;

			10100: dout = 12'h000;
			10101: dout = 12'h000;
			10102: dout = 12'h000;
			10103: dout = 12'h000;
			10104: dout = 12'h000;
			10105: dout = 12'h000;
			10106: dout = 12'h000;
			10107: dout = 12'h000;
			10108: dout = 12'h000;
			10109: dout = 12'h000;
			10110: dout = 12'h000;
			10111: dout = 12'h000;
			10112: dout = 12'h000;
			10113: dout = 12'h000;
			10114: dout = 12'h000;
			10115: dout = 12'h000;
			10116: dout = 12'h000;
			10117: dout = 12'h000;

			10118: dout = 12'h000;
			10119: dout = 12'h000;
			10120: dout = 12'h000;
			10121: dout = 12'h000;
			10122: dout = 12'h000;
			10123: dout = 12'h114;
			10124: dout = 12'h34c;
			10125: dout = 12'h114;
			10126: dout = 12'h000;
			10127: dout = 12'h113;
			10128: dout = 12'h34c;
			10129: dout = 12'h34c;
			10130: dout = 12'h238;
			10131: dout = 12'h002;
			10132: dout = 12'h000;
			10133: dout = 12'h000;
			10134: dout = 12'h000;
			10135: dout = 12'h000;

			10136: dout = 12'h000;
			10137: dout = 12'h000;
			10138: dout = 12'h000;
			10139: dout = 12'h000;
			10140: dout = 12'h115;
			10141: dout = 12'h34a;
			10142: dout = 12'h35a;
			10143: dout = 12'h000;
			10144: dout = 12'h000;
			10145: dout = 12'h258;
			10146: dout = 12'h34a;
			10147: dout = 12'h226;
			10148: dout = 12'h001;
			10149: dout = 12'h237;
			10150: dout = 12'h114;
			10151: dout = 12'h000;
			10152: dout = 12'h000;
			10153: dout = 12'h000;

			10154: dout = 12'h000;
			10155: dout = 12'h000;
			10156: dout = 12'h000;
			10157: dout = 12'h000;
			10158: dout = 12'h237;
			10159: dout = 12'h46e;
			10160: dout = 12'h36a;
			10161: dout = 12'h000;
			10162: dout = 12'h000;
			10163: dout = 12'h36b;
			10164: dout = 12'h011;
			10165: dout = 12'h000;
			10166: dout = 12'h000;
			10167: dout = 12'h238;
			10168: dout = 12'h34a;
			10169: dout = 12'h113;
			10170: dout = 12'h001;
			10171: dout = 12'h000;

			10172: dout = 12'h000;
			10173: dout = 12'h000;
			10174: dout = 12'h000;
			10175: dout = 12'h000;
			10176: dout = 12'h000;
			10177: dout = 12'h000;
			10178: dout = 12'h248;
			10179: dout = 12'h000;
			10180: dout = 12'h000;
			10181: dout = 12'h000;
			10182: dout = 12'h000;
			10183: dout = 12'h000;
			10184: dout = 12'h000;
			10185: dout = 12'h000;
			10186: dout = 12'h000;
			10187: dout = 12'h229;
			10188: dout = 12'h002;
			10189: dout = 12'h000;

			10190: dout = 12'h000;
			10191: dout = 12'h000;
			10192: dout = 12'h000;
			10193: dout = 12'h000;
			10194: dout = 12'h000;
			10195: dout = 12'h000;
			10196: dout = 12'h000;
			10197: dout = 12'h000;
			10198: dout = 12'h000;
			10199: dout = 12'h000;
			10200: dout = 12'h000;
			10201: dout = 12'h000;
			10202: dout = 12'h000;
			10203: dout = 12'h123;
			10204: dout = 12'h247;
			10205: dout = 12'h000;
			10206: dout = 12'h000;
			10207: dout = 12'h001;

			10208: dout = 12'h000;
			10209: dout = 12'h000;
			10210: dout = 12'h000;
			10211: dout = 12'h000;
			10212: dout = 12'h000;
			10213: dout = 12'h000;
			10214: dout = 12'h000;
			10215: dout = 12'h000;
			10216: dout = 12'h000;
			10217: dout = 12'h000;
			10218: dout = 12'h000;
			10219: dout = 12'h000;
			10220: dout = 12'h000;
			10221: dout = 12'h247;
			10222: dout = 12'h48e;
			10223: dout = 12'h248;
			10224: dout = 12'h000;
			10225: dout = 12'h000;

			10226: dout = 12'h000;
			10227: dout = 12'h000;
			10228: dout = 12'h000;
			10229: dout = 12'h000;
			10230: dout = 12'h000;
			10231: dout = 12'h000;
			10232: dout = 12'h000;
			10233: dout = 12'h000;
			10234: dout = 12'h000;
			10235: dout = 12'h000;
			10236: dout = 12'h000;
			10237: dout = 12'h000;
			10238: dout = 12'h000;
			10239: dout = 12'h000;
			10240: dout = 12'h000;
			10241: dout = 12'h000;
			10242: dout = 12'h000;
			10243: dout = 12'h000;

			10244: dout = 12'h000;
			10245: dout = 12'h012;
			10246: dout = 12'h226;
			10247: dout = 12'h237;
			10248: dout = 12'h123;
			10249: dout = 12'h000;
			10250: dout = 12'h000;
			10251: dout = 12'h000;
			10252: dout = 12'h000;
			10253: dout = 12'h000;
			10254: dout = 12'h000;
			10255: dout = 12'h000;
			10256: dout = 12'h000;
			10257: dout = 12'h000;
			10258: dout = 12'h000;
			10259: dout = 12'h247;
			10260: dout = 12'h226;
			10261: dout = 12'h001;

			10262: dout = 12'h000;
			10263: dout = 12'h113;
			10264: dout = 12'h34b;
			10265: dout = 12'h47d;
			10266: dout = 12'h247;
			10267: dout = 12'h000;
			10268: dout = 12'h000;
			10269: dout = 12'h000;
			10270: dout = 12'h000;
			10271: dout = 12'h000;
			10272: dout = 12'h000;
			10273: dout = 12'h000;
			10274: dout = 12'h000;
			10275: dout = 12'h000;
			10276: dout = 12'h000;
			10277: dout = 12'h48e;
			10278: dout = 12'h45d;
			10279: dout = 12'h113;

			10280: dout = 12'h000;
			10281: dout = 12'h002;
			10282: dout = 12'h228;
			10283: dout = 12'h237;
			10284: dout = 12'h000;
			10285: dout = 12'h000;
			10286: dout = 12'h000;
			10287: dout = 12'h000;
			10288: dout = 12'h000;
			10289: dout = 12'h000;
			10290: dout = 12'h000;
			10291: dout = 12'h000;
			10292: dout = 12'h000;
			10293: dout = 12'h000;
			10294: dout = 12'h000;
			10295: dout = 12'h113;
			10296: dout = 12'h34b;
			10297: dout = 12'h002;

			10298: dout = 12'h000;
			10299: dout = 12'h000;
			10300: dout = 12'h000;
			10301: dout = 12'h000;
			10302: dout = 12'h000;
			10303: dout = 12'h000;
			10304: dout = 12'h000;
			10305: dout = 12'h000;
			10306: dout = 12'h000;
			10307: dout = 12'h000;
			10308: dout = 12'h000;
			10309: dout = 12'h000;
			10310: dout = 12'h000;
			10311: dout = 12'h000;
			10312: dout = 12'h000;
			10313: dout = 12'h001;
			10314: dout = 12'h113;
			10315: dout = 12'h000;

			10316: dout = 12'h000;
			10317: dout = 12'h000;
			10318: dout = 12'h000;
			10319: dout = 12'h000;
			10320: dout = 12'h000;
			10321: dout = 12'h000;
			10322: dout = 12'h000;
			10323: dout = 12'h000;
			10324: dout = 12'h000;
			10325: dout = 12'h000;
			10326: dout = 12'h000;
			10327: dout = 12'h000;
			10328: dout = 12'h000;
			10329: dout = 12'h000;
			10330: dout = 12'h000;
			10331: dout = 12'h000;
			10332: dout = 12'h000;
			10333: dout = 12'h000;

			10334: dout = 12'h000;
			10335: dout = 12'h000;
			10336: dout = 12'h000;
			10337: dout = 12'h000;
			10338: dout = 12'h000;
			10339: dout = 12'h000;
			10340: dout = 12'h000;
			10341: dout = 12'h000;
			10342: dout = 12'h000;
			10343: dout = 12'h000;
			10344: dout = 12'h000;
			10345: dout = 12'h000;
			10346: dout = 12'h000;
			10347: dout = 12'h000;
			10348: dout = 12'h000;
			10349: dout = 12'h000;
			10350: dout = 12'h000;
			10351: dout = 12'h000;

			10352: dout = 12'h000;
			10353: dout = 12'h000;
			10354: dout = 12'h000;
			10355: dout = 12'h000;
			10356: dout = 12'h000;
			10357: dout = 12'h000;
			10358: dout = 12'h000;
			10359: dout = 12'h000;
			10360: dout = 12'h000;
			10361: dout = 12'h000;
			10362: dout = 12'h000;
			10363: dout = 12'h000;
			10364: dout = 12'h000;
			10365: dout = 12'h000;
			10366: dout = 12'h000;
			10367: dout = 12'h000;
			10368: dout = 12'h000;
			10369: dout = 12'h000;

			10370: dout = 12'h000;
			10371: dout = 12'h000;
			10372: dout = 12'h000;
			10373: dout = 12'h000;
			10374: dout = 12'h000;
			10375: dout = 12'h000;
			10376: dout = 12'h000;
			10377: dout = 12'h000;
			10378: dout = 12'h000;
			10379: dout = 12'h000;
			10380: dout = 12'h000;
			10381: dout = 12'h000;
			10382: dout = 12'h000;
			10383: dout = 12'h000;
			10384: dout = 12'h000;
			10385: dout = 12'h000;
			10386: dout = 12'h000;
			10387: dout = 12'h000;

			10388: dout = 12'h000;
			10389: dout = 12'h115;
			10390: dout = 12'h35c;
			10391: dout = 12'h36b;
			10392: dout = 12'h001;
			10393: dout = 12'h000;
			10394: dout = 12'h000;
			10395: dout = 12'h000;
			10396: dout = 12'h000;
			10397: dout = 12'h000;
			10398: dout = 12'h000;
			10399: dout = 12'h000;
			10400: dout = 12'h000;
			10401: dout = 12'h011;
			10402: dout = 12'h36b;
			10403: dout = 12'h36b;
			10404: dout = 12'h000;
			10405: dout = 12'h000;

			10406: dout = 12'h000;
			10407: dout = 12'h000;
			10408: dout = 12'h114;
			10409: dout = 12'h33b;
			10410: dout = 12'h113;
			10411: dout = 12'h000;
			10412: dout = 12'h011;
			10413: dout = 12'h123;
			10414: dout = 12'h000;
			10415: dout = 12'h000;
			10416: dout = 12'h000;
			10417: dout = 12'h000;
			10418: dout = 12'h135;
			10419: dout = 12'h123;
			10420: dout = 12'h35b;
			10421: dout = 12'h33a;
			10422: dout = 12'h002;
			10423: dout = 12'h000;

			10424: dout = 12'h000;
			10425: dout = 12'h000;
			10426: dout = 12'h001;
			10427: dout = 12'h002;
			10428: dout = 12'h000;
			10429: dout = 12'h000;
			10430: dout = 12'h37b;
			10431: dout = 12'h47c;
			10432: dout = 12'h012;
			10433: dout = 12'h000;
			10434: dout = 12'h000;
			10435: dout = 12'h248;
			10436: dout = 12'h47d;
			10437: dout = 12'h125;
			10438: dout = 12'h125;
			10439: dout = 12'h002;
			10440: dout = 12'h000;
			10441: dout = 12'h000;

			10442: dout = 12'h000;
			10443: dout = 12'h000;
			10444: dout = 12'h000;
			10445: dout = 12'h000;
			10446: dout = 12'h001;
			10447: dout = 12'h237;
			10448: dout = 12'h46e;
			10449: dout = 12'h47e;
			10450: dout = 12'h123;
			10451: dout = 12'h000;
			10452: dout = 12'h000;
			10453: dout = 12'h35a;
			10454: dout = 12'h45d;
			10455: dout = 12'h124;
			10456: dout = 12'h002;
			10457: dout = 12'h000;
			10458: dout = 12'h000;
			10459: dout = 12'h000;

			10460: dout = 12'h000;
			10461: dout = 12'h000;
			10462: dout = 12'h000;
			10463: dout = 12'h000;
			10464: dout = 12'h000;
			10465: dout = 12'h013;
			10466: dout = 12'h239;
			10467: dout = 12'h249;
			10468: dout = 12'h011;
			10469: dout = 12'h000;
			10470: dout = 12'h113;
			10471: dout = 12'h34a;
			10472: dout = 12'h227;
			10473: dout = 12'h002;
			10474: dout = 12'h000;
			10475: dout = 12'h000;
			10476: dout = 12'h000;
			10477: dout = 12'h000;

			10478: dout = 12'h000;
			10479: dout = 12'h000;
			10480: dout = 12'h000;
			10481: dout = 12'h000;
			10482: dout = 12'h000;
			10483: dout = 12'h000;
			10484: dout = 12'h001;
			10485: dout = 12'h001;
			10486: dout = 12'h000;
			10487: dout = 12'h000;
			10488: dout = 12'h001;
			10489: dout = 12'h126;
			10490: dout = 12'h000;
			10491: dout = 12'h000;
			10492: dout = 12'h000;
			10493: dout = 12'h000;
			10494: dout = 12'h000;
			10495: dout = 12'h000;

			10496: dout = 12'h000;
			10497: dout = 12'h000;
			10498: dout = 12'h000;
			10499: dout = 12'h000;
			10500: dout = 12'h000;
			10501: dout = 12'h000;
			10502: dout = 12'h000;
			10503: dout = 12'h000;
			10504: dout = 12'h000;
			10505: dout = 12'h001;
			10506: dout = 12'h113;
			10507: dout = 12'h000;
			10508: dout = 12'h000;
			10509: dout = 12'h000;
			10510: dout = 12'h000;
			10511: dout = 12'h000;
			10512: dout = 12'h000;
			10513: dout = 12'h000;

			10514: dout = 12'h000;
			10515: dout = 12'h000;
			10516: dout = 12'h000;
			10517: dout = 12'h000;
			10518: dout = 12'h000;
			10519: dout = 12'h000;
			10520: dout = 12'h000;
			10521: dout = 12'h000;
			10522: dout = 12'h000;
			10523: dout = 12'h000;
			10524: dout = 12'h001;
			10525: dout = 12'h000;
			10526: dout = 12'h000;
			10527: dout = 12'h000;
			10528: dout = 12'h000;
			10529: dout = 12'h000;
			10530: dout = 12'h000;
			10531: dout = 12'h000;

			10532: dout = 12'h000;
			10533: dout = 12'h000;
			10534: dout = 12'h000;
			10535: dout = 12'h000;
			10536: dout = 12'h000;
			10537: dout = 12'h000;
			10538: dout = 12'h000;
			10539: dout = 12'h000;
			10540: dout = 12'h000;
			10541: dout = 12'h000;
			10542: dout = 12'h000;
			10543: dout = 12'h000;
			10544: dout = 12'h000;
			10545: dout = 12'h000;
			10546: dout = 12'h000;
			10547: dout = 12'h000;
			10548: dout = 12'h000;
			10549: dout = 12'h000;

			10550: dout = 12'h000;
			10551: dout = 12'h000;
			10552: dout = 12'h000;
			10553: dout = 12'h000;
			10554: dout = 12'h000;
			10555: dout = 12'h000;
			10556: dout = 12'h000;
			10557: dout = 12'h000;
			10558: dout = 12'h000;
			10559: dout = 12'h000;
			10560: dout = 12'h000;
			10561: dout = 12'h000;
			10562: dout = 12'h000;
			10563: dout = 12'h000;
			10564: dout = 12'h000;
			10565: dout = 12'h000;
			10566: dout = 12'h000;
			10567: dout = 12'h000;
			10568: dout = 12'h000;
			10569: dout = 12'h000;
			10570: dout = 12'h000;
			10571: dout = 12'h000;
			10572: dout = 12'h000;
			10573: dout = 12'h000;
			10574: dout = 12'h000;
			10575: dout = 12'h000;
			10576: dout = 12'h000;
			10577: dout = 12'h000;
			10578: dout = 12'h000;
			10579: dout = 12'h000;
			10580: dout = 12'h000;
			10581: dout = 12'h000;
			10582: dout = 12'h000;
			10583: dout = 12'h000;
			10584: dout = 12'h000;
			10585: dout = 12'h000;
			10586: dout = 12'h000;
			10587: dout = 12'h000;
			10588: dout = 12'h000;
			10589: dout = 12'h000;
			10590: dout = 12'h000;
			10591: dout = 12'h000;
			10592: dout = 12'h000;
			10593: dout = 12'h000;
			10594: dout = 12'h000;
			10595: dout = 12'h000;
			10596: dout = 12'h000;
			10597: dout = 12'h000;
			10598: dout = 12'h000;
			10599: dout = 12'h000;

			10600: dout = 12'h000;
			10601: dout = 12'h000;
			10602: dout = 12'h000;
			10603: dout = 12'h000;
			10604: dout = 12'h000;
			10605: dout = 12'h000;
			10606: dout = 12'h000;
			10607: dout = 12'h000;
			10608: dout = 12'h000;
			10609: dout = 12'h000;
			10610: dout = 12'h000;
			10611: dout = 12'h000;
			10612: dout = 12'h000;
			10613: dout = 12'h000;
			10614: dout = 12'h000;
			10615: dout = 12'h000;
			10616: dout = 12'h000;
			10617: dout = 12'h000;
			10618: dout = 12'h000;
			10619: dout = 12'h000;
			10620: dout = 12'h000;
			10621: dout = 12'h000;
			10622: dout = 12'h000;
			10623: dout = 12'h000;
			10624: dout = 12'h000;
			10625: dout = 12'h000;
			10626: dout = 12'h000;
			10627: dout = 12'h000;
			10628: dout = 12'h000;
			10629: dout = 12'h000;
			10630: dout = 12'h000;
			10631: dout = 12'h000;
			10632: dout = 12'h000;
			10633: dout = 12'h000;
			10634: dout = 12'h000;
			10635: dout = 12'h000;
			10636: dout = 12'h000;
			10637: dout = 12'h000;
			10638: dout = 12'h000;
			10639: dout = 12'h000;
			10640: dout = 12'h000;
			10641: dout = 12'h000;
			10642: dout = 12'h000;
			10643: dout = 12'h000;
			10644: dout = 12'h000;
			10645: dout = 12'h000;
			10646: dout = 12'h000;
			10647: dout = 12'h000;
			10648: dout = 12'h000;
			10649: dout = 12'h000;

			10650: dout = 12'h000;
			10651: dout = 12'h000;
			10652: dout = 12'h000;
			10653: dout = 12'h000;
			10654: dout = 12'h000;
			10655: dout = 12'h000;
			10656: dout = 12'h000;
			10657: dout = 12'h000;
			10658: dout = 12'h000;
			10659: dout = 12'h000;
			10660: dout = 12'h000;
			10661: dout = 12'h000;
			10662: dout = 12'h000;
			10663: dout = 12'h000;
			10664: dout = 12'h000;
			10665: dout = 12'h000;
			10666: dout = 12'h000;
			10667: dout = 12'h000;
			10668: dout = 12'h000;
			10669: dout = 12'h000;
			10670: dout = 12'h000;
			10671: dout = 12'h000;
			10672: dout = 12'h000;
			10673: dout = 12'h000;
			10674: dout = 12'h000;
			10675: dout = 12'h000;
			10676: dout = 12'h000;
			10677: dout = 12'h000;
			10678: dout = 12'h000;
			10679: dout = 12'h000;
			10680: dout = 12'h000;
			10681: dout = 12'h000;
			10682: dout = 12'h000;
			10683: dout = 12'h000;
			10684: dout = 12'h000;
			10685: dout = 12'h000;
			10686: dout = 12'h000;
			10687: dout = 12'h000;
			10688: dout = 12'h000;
			10689: dout = 12'h000;
			10690: dout = 12'h000;
			10691: dout = 12'h000;
			10692: dout = 12'h000;
			10693: dout = 12'h000;
			10694: dout = 12'h000;
			10695: dout = 12'h000;
			10696: dout = 12'h000;
			10697: dout = 12'h000;
			10698: dout = 12'h000;
			10699: dout = 12'h000;

			10700: dout = 12'h000;
			10701: dout = 12'h000;
			10702: dout = 12'h000;
			10703: dout = 12'h000;
			10704: dout = 12'h000;
			10705: dout = 12'h000;
			10706: dout = 12'h000;
			10707: dout = 12'h000;
			10708: dout = 12'h000;
			10709: dout = 12'h000;
			10710: dout = 12'h000;
			10711: dout = 12'h000;
			10712: dout = 12'h000;
			10713: dout = 12'h000;
			10714: dout = 12'h000;
			10715: dout = 12'h000;
			10716: dout = 12'h000;
			10717: dout = 12'h000;
			10718: dout = 12'h000;
			10719: dout = 12'h000;
			10720: dout = 12'h000;
			10721: dout = 12'h000;
			10722: dout = 12'h000;
			10723: dout = 12'h000;
			10724: dout = 12'h000;
			10725: dout = 12'h000;
			10726: dout = 12'h000;
			10727: dout = 12'h000;
			10728: dout = 12'h000;
			10729: dout = 12'h000;
			10730: dout = 12'h000;
			10731: dout = 12'h000;
			10732: dout = 12'h000;
			10733: dout = 12'h000;
			10734: dout = 12'h000;
			10735: dout = 12'h000;
			10736: dout = 12'h000;
			10737: dout = 12'h000;
			10738: dout = 12'h000;
			10739: dout = 12'h000;
			10740: dout = 12'h000;
			10741: dout = 12'h000;
			10742: dout = 12'h000;
			10743: dout = 12'h000;
			10744: dout = 12'h000;
			10745: dout = 12'h000;
			10746: dout = 12'h000;
			10747: dout = 12'h000;
			10748: dout = 12'h000;
			10749: dout = 12'h000;

			10750: dout = 12'h000;
			10751: dout = 12'h000;
			10752: dout = 12'h000;
			10753: dout = 12'h000;
			10754: dout = 12'h000;
			10755: dout = 12'h000;
			10756: dout = 12'h000;
			10757: dout = 12'h000;
			10758: dout = 12'h000;
			10759: dout = 12'h000;
			10760: dout = 12'h000;
			10761: dout = 12'h000;
			10762: dout = 12'h000;
			10763: dout = 12'h000;
			10764: dout = 12'h000;
			10765: dout = 12'h000;
			10766: dout = 12'h000;
			10767: dout = 12'h000;
			10768: dout = 12'h000;
			10769: dout = 12'h000;
			10770: dout = 12'h000;
			10771: dout = 12'h000;
			10772: dout = 12'h000;
			10773: dout = 12'h000;
			10774: dout = 12'h000;
			10775: dout = 12'h000;
			10776: dout = 12'h000;
			10777: dout = 12'h000;
			10778: dout = 12'h000;
			10779: dout = 12'h000;
			10780: dout = 12'h000;
			10781: dout = 12'h000;
			10782: dout = 12'h000;
			10783: dout = 12'h000;
			10784: dout = 12'h000;
			10785: dout = 12'h000;
			10786: dout = 12'h000;
			10787: dout = 12'h000;
			10788: dout = 12'h000;
			10789: dout = 12'h000;
			10790: dout = 12'h000;
			10791: dout = 12'h000;
			10792: dout = 12'h000;
			10793: dout = 12'h000;
			10794: dout = 12'h000;
			10795: dout = 12'h000;
			10796: dout = 12'h000;
			10797: dout = 12'h000;
			10798: dout = 12'h000;
			10799: dout = 12'h000;

			10800: dout = 12'h000;
			10801: dout = 12'h000;
			10802: dout = 12'h000;
			10803: dout = 12'h000;
			10804: dout = 12'h000;
			10805: dout = 12'h000;
			10806: dout = 12'h000;
			10807: dout = 12'h000;
			10808: dout = 12'h000;
			10809: dout = 12'h000;
			10810: dout = 12'h000;
			10811: dout = 12'h000;
			10812: dout = 12'h000;
			10813: dout = 12'h000;
			10814: dout = 12'h000;
			10815: dout = 12'h000;
			10816: dout = 12'h000;
			10817: dout = 12'h000;
			10818: dout = 12'h000;
			10819: dout = 12'h000;
			10820: dout = 12'h000;
			10821: dout = 12'h000;
			10822: dout = 12'h000;
			10823: dout = 12'h000;
			10824: dout = 12'h000;
			10825: dout = 12'h000;
			10826: dout = 12'h000;
			10827: dout = 12'h000;
			10828: dout = 12'h000;
			10829: dout = 12'h000;
			10830: dout = 12'h000;
			10831: dout = 12'h000;
			10832: dout = 12'h000;
			10833: dout = 12'h000;
			10834: dout = 12'h000;
			10835: dout = 12'h000;
			10836: dout = 12'h000;
			10837: dout = 12'h000;
			10838: dout = 12'h000;
			10839: dout = 12'h000;
			10840: dout = 12'h000;
			10841: dout = 12'h000;
			10842: dout = 12'h000;
			10843: dout = 12'h000;
			10844: dout = 12'h000;
			10845: dout = 12'h000;
			10846: dout = 12'h000;
			10847: dout = 12'h000;
			10848: dout = 12'h000;
			10849: dout = 12'h000;

			10850: dout = 12'h000;
			10851: dout = 12'h000;
			10852: dout = 12'h000;
			10853: dout = 12'h000;
			10854: dout = 12'h000;
			10855: dout = 12'h000;
			10856: dout = 12'h000;
			10857: dout = 12'h000;
			10858: dout = 12'h000;
			10859: dout = 12'h000;
			10860: dout = 12'h000;
			10861: dout = 12'h000;
			10862: dout = 12'h000;
			10863: dout = 12'h000;
			10864: dout = 12'h000;
			10865: dout = 12'h000;
			10866: dout = 12'h000;
			10867: dout = 12'h000;
			10868: dout = 12'h000;
			10869: dout = 12'h000;
			10870: dout = 12'h000;
			10871: dout = 12'h000;
			10872: dout = 12'h000;
			10873: dout = 12'h000;
			10874: dout = 12'h000;
			10875: dout = 12'h000;
			10876: dout = 12'h000;
			10877: dout = 12'h000;
			10878: dout = 12'h000;
			10879: dout = 12'h000;
			10880: dout = 12'h000;
			10881: dout = 12'h000;
			10882: dout = 12'h000;
			10883: dout = 12'h000;
			10884: dout = 12'h000;
			10885: dout = 12'h000;
			10886: dout = 12'h000;
			10887: dout = 12'h000;
			10888: dout = 12'h000;
			10889: dout = 12'h000;
			10890: dout = 12'h000;
			10891: dout = 12'h000;
			10892: dout = 12'h000;
			10893: dout = 12'h000;
			10894: dout = 12'h000;
			10895: dout = 12'h000;
			10896: dout = 12'h000;
			10897: dout = 12'h000;
			10898: dout = 12'h000;
			10899: dout = 12'h000;

			10900: dout = 12'h000;
			10901: dout = 12'h000;
			10902: dout = 12'h000;
			10903: dout = 12'h000;
			10904: dout = 12'h000;
			10905: dout = 12'h000;
			10906: dout = 12'h000;
			10907: dout = 12'h000;
			10908: dout = 12'h000;
			10909: dout = 12'h000;
			10910: dout = 12'h000;
			10911: dout = 12'h000;
			10912: dout = 12'h000;
			10913: dout = 12'h000;
			10914: dout = 12'h000;
			10915: dout = 12'h000;
			10916: dout = 12'h000;
			10917: dout = 12'h000;
			10918: dout = 12'h000;
			10919: dout = 12'h000;
			10920: dout = 12'h000;
			10921: dout = 12'h000;
			10922: dout = 12'h000;
			10923: dout = 12'h000;
			10924: dout = 12'h000;
			10925: dout = 12'h000;
			10926: dout = 12'h000;
			10927: dout = 12'h000;
			10928: dout = 12'h000;
			10929: dout = 12'h000;
			10930: dout = 12'h000;
			10931: dout = 12'h000;
			10932: dout = 12'h000;
			10933: dout = 12'h000;
			10934: dout = 12'h000;
			10935: dout = 12'h000;
			10936: dout = 12'h000;
			10937: dout = 12'h000;
			10938: dout = 12'h000;
			10939: dout = 12'h000;
			10940: dout = 12'h000;
			10941: dout = 12'h000;
			10942: dout = 12'h000;
			10943: dout = 12'h000;
			10944: dout = 12'h000;
			10945: dout = 12'h000;
			10946: dout = 12'h000;
			10947: dout = 12'h000;
			10948: dout = 12'h000;
			10949: dout = 12'h000;

			10950: dout = 12'h000;
			10951: dout = 12'h000;
			10952: dout = 12'h000;
			10953: dout = 12'h000;
			10954: dout = 12'h000;
			10955: dout = 12'h000;
			10956: dout = 12'h000;
			10957: dout = 12'h000;
			10958: dout = 12'h000;
			10959: dout = 12'h000;
			10960: dout = 12'h000;
			10961: dout = 12'h000;
			10962: dout = 12'h000;
			10963: dout = 12'h000;
			10964: dout = 12'h000;
			10965: dout = 12'h000;
			10966: dout = 12'h000;
			10967: dout = 12'h000;
			10968: dout = 12'h000;
			10969: dout = 12'h000;
			10970: dout = 12'h000;
			10971: dout = 12'h000;
			10972: dout = 12'h000;
			10973: dout = 12'h000;
			10974: dout = 12'h000;
			10975: dout = 12'h000;
			10976: dout = 12'h000;
			10977: dout = 12'h000;
			10978: dout = 12'h000;
			10979: dout = 12'h000;
			10980: dout = 12'h000;
			10981: dout = 12'h000;
			10982: dout = 12'h000;
			10983: dout = 12'h000;
			10984: dout = 12'h000;
			10985: dout = 12'h000;
			10986: dout = 12'h000;
			10987: dout = 12'h000;
			10988: dout = 12'h000;
			10989: dout = 12'h000;
			10990: dout = 12'h000;
			10991: dout = 12'h000;
			10992: dout = 12'h000;
			10993: dout = 12'h000;
			10994: dout = 12'h000;
			10995: dout = 12'h000;
			10996: dout = 12'h000;
			10997: dout = 12'h000;
			10998: dout = 12'h000;
			10999: dout = 12'h000;

			11000: dout = 12'h000;
			11001: dout = 12'h000;
			11002: dout = 12'h000;
			11003: dout = 12'h000;
			11004: dout = 12'h000;
			11005: dout = 12'h000;
			11006: dout = 12'h000;
			11007: dout = 12'h000;
			11008: dout = 12'h000;
			11009: dout = 12'h000;
			11010: dout = 12'h000;
			11011: dout = 12'h000;
			11012: dout = 12'h000;
			11013: dout = 12'h000;
			11014: dout = 12'h000;
			11015: dout = 12'h000;
			11016: dout = 12'h000;
			11017: dout = 12'h000;
			11018: dout = 12'h000;
			11019: dout = 12'h000;
			11020: dout = 12'h000;
			11021: dout = 12'h000;
			11022: dout = 12'h000;
			11023: dout = 12'h000;
			11024: dout = 12'h000;
			11025: dout = 12'h000;
			11026: dout = 12'h000;
			11027: dout = 12'h000;
			11028: dout = 12'h000;
			11029: dout = 12'h000;
			11030: dout = 12'h000;
			11031: dout = 12'h000;
			11032: dout = 12'h000;
			11033: dout = 12'h000;
			11034: dout = 12'h000;
			11035: dout = 12'h000;
			11036: dout = 12'h000;
			11037: dout = 12'h000;
			11038: dout = 12'h000;
			11039: dout = 12'h000;
			11040: dout = 12'h000;
			11041: dout = 12'h000;
			11042: dout = 12'h000;
			11043: dout = 12'h000;
			11044: dout = 12'h000;
			11045: dout = 12'h000;
			11046: dout = 12'h000;
			11047: dout = 12'h000;
			11048: dout = 12'h000;
			11049: dout = 12'h000;

			11050: dout = 12'h000;
			11051: dout = 12'h000;
			11052: dout = 12'h000;
			11053: dout = 12'h000;
			11054: dout = 12'h000;
			11055: dout = 12'h000;
			11056: dout = 12'h000;
			11057: dout = 12'h000;
			11058: dout = 12'h000;
			11059: dout = 12'h000;
			11060: dout = 12'h000;
			11061: dout = 12'h000;
			11062: dout = 12'h000;
			11063: dout = 12'h000;
			11064: dout = 12'h000;
			11065: dout = 12'h000;
			11066: dout = 12'h000;
			11067: dout = 12'h000;
			11068: dout = 12'h000;
			11069: dout = 12'h000;
			11070: dout = 12'h000;
			11071: dout = 12'h000;
			11072: dout = 12'h000;
			11073: dout = 12'h000;
			11074: dout = 12'h000;
			11075: dout = 12'h000;
			11076: dout = 12'h555;
			11077: dout = 12'h333;
			11078: dout = 12'h000;
			11079: dout = 12'h000;
			11080: dout = 12'h000;
			11081: dout = 12'h000;
			11082: dout = 12'h000;
			11083: dout = 12'h000;
			11084: dout = 12'h000;
			11085: dout = 12'h000;
			11086: dout = 12'h000;
			11087: dout = 12'h000;
			11088: dout = 12'h000;
			11089: dout = 12'h000;
			11090: dout = 12'h000;
			11091: dout = 12'h000;
			11092: dout = 12'h000;
			11093: dout = 12'h000;
			11094: dout = 12'h000;
			11095: dout = 12'h000;
			11096: dout = 12'h000;
			11097: dout = 12'h000;
			11098: dout = 12'h000;
			11099: dout = 12'h000;

			11100: dout = 12'h000;
			11101: dout = 12'h000;
			11102: dout = 12'h000;
			11103: dout = 12'h000;
			11104: dout = 12'h000;
			11105: dout = 12'h000;
			11106: dout = 12'h000;
			11107: dout = 12'h000;
			11108: dout = 12'h000;
			11109: dout = 12'h000;
			11110: dout = 12'h000;
			11111: dout = 12'h000;
			11112: dout = 12'h000;
			11113: dout = 12'h000;
			11114: dout = 12'h000;
			11115: dout = 12'h000;
			11116: dout = 12'h000;
			11117: dout = 12'h000;
			11118: dout = 12'h000;
			11119: dout = 12'h000;
			11120: dout = 12'h000;
			11121: dout = 12'h000;
			11122: dout = 12'h000;
			11123: dout = 12'h000;
			11124: dout = 12'h000;
			11125: dout = 12'hbbb;
			11126: dout = 12'hfff;
			11127: dout = 12'hfff;
			11128: dout = 12'h444;
			11129: dout = 12'h000;
			11130: dout = 12'h000;
			11131: dout = 12'h000;
			11132: dout = 12'h000;
			11133: dout = 12'h000;
			11134: dout = 12'h000;
			11135: dout = 12'h000;
			11136: dout = 12'h000;
			11137: dout = 12'h000;
			11138: dout = 12'h000;
			11139: dout = 12'h000;
			11140: dout = 12'h000;
			11141: dout = 12'h000;
			11142: dout = 12'h000;
			11143: dout = 12'h000;
			11144: dout = 12'h000;
			11145: dout = 12'h000;
			11146: dout = 12'h000;
			11147: dout = 12'h000;
			11148: dout = 12'h000;
			11149: dout = 12'h000;

			11150: dout = 12'h000;
			11151: dout = 12'h000;
			11152: dout = 12'h000;
			11153: dout = 12'h000;
			11154: dout = 12'h000;
			11155: dout = 12'h000;
			11156: dout = 12'h000;
			11157: dout = 12'h000;
			11158: dout = 12'h000;
			11159: dout = 12'h000;
			11160: dout = 12'h000;
			11161: dout = 12'h000;
			11162: dout = 12'h000;
			11163: dout = 12'h000;
			11164: dout = 12'h000;
			11165: dout = 12'h000;
			11166: dout = 12'h000;
			11167: dout = 12'h000;
			11168: dout = 12'h000;
			11169: dout = 12'h000;
			11170: dout = 12'h000;
			11171: dout = 12'h000;
			11172: dout = 12'h000;
			11173: dout = 12'h000;
			11174: dout = 12'h000;
			11175: dout = 12'hfff;
			11176: dout = 12'h776;
			11177: dout = 12'hfff;
			11178: dout = 12'h666;
			11179: dout = 12'h000;
			11180: dout = 12'h000;
			11181: dout = 12'h000;
			11182: dout = 12'h000;
			11183: dout = 12'h000;
			11184: dout = 12'h000;
			11185: dout = 12'h000;
			11186: dout = 12'h000;
			11187: dout = 12'h000;
			11188: dout = 12'h000;
			11189: dout = 12'h000;
			11190: dout = 12'h000;
			11191: dout = 12'h000;
			11192: dout = 12'h000;
			11193: dout = 12'h000;
			11194: dout = 12'h000;
			11195: dout = 12'h000;
			11196: dout = 12'h000;
			11197: dout = 12'h000;
			11198: dout = 12'h000;
			11199: dout = 12'h000;

			11200: dout = 12'h000;
			11201: dout = 12'h000;
			11202: dout = 12'h000;
			11203: dout = 12'h000;
			11204: dout = 12'h000;
			11205: dout = 12'h000;
			11206: dout = 12'h000;
			11207: dout = 12'h000;
			11208: dout = 12'h000;
			11209: dout = 12'h000;
			11210: dout = 12'h000;
			11211: dout = 12'h000;
			11212: dout = 12'h000;
			11213: dout = 12'h000;
			11214: dout = 12'h000;
			11215: dout = 12'h000;
			11216: dout = 12'h000;
			11217: dout = 12'h000;
			11218: dout = 12'hbbc;
			11219: dout = 12'hddd;
			11220: dout = 12'h111;
			11221: dout = 12'h000;
			11222: dout = 12'h000;
			11223: dout = 12'h000;
			11224: dout = 12'h222;
			11225: dout = 12'hfff;
			11226: dout = 12'h211;
			11227: dout = 12'hfff;
			11228: dout = 12'h666;
			11229: dout = 12'h000;
			11230: dout = 12'h000;
			11231: dout = 12'h000;
			11232: dout = 12'h000;
			11233: dout = 12'h000;
			11234: dout = 12'h888;
			11235: dout = 12'heee;
			11236: dout = 12'h777;
			11237: dout = 12'h000;
			11238: dout = 12'h000;
			11239: dout = 12'h000;
			11240: dout = 12'h000;
			11241: dout = 12'h000;
			11242: dout = 12'h000;
			11243: dout = 12'h000;
			11244: dout = 12'h000;
			11245: dout = 12'h000;
			11246: dout = 12'h000;
			11247: dout = 12'h000;
			11248: dout = 12'h000;
			11249: dout = 12'h000;

			11250: dout = 12'h000;
			11251: dout = 12'h000;
			11252: dout = 12'h000;
			11253: dout = 12'h000;
			11254: dout = 12'h000;
			11255: dout = 12'h000;
			11256: dout = 12'h000;
			11257: dout = 12'h000;
			11258: dout = 12'h000;
			11259: dout = 12'h000;
			11260: dout = 12'h000;
			11261: dout = 12'h000;
			11262: dout = 12'h000;
			11263: dout = 12'hddd;
			11264: dout = 12'heee;
			11265: dout = 12'h000;
			11266: dout = 12'h000;
			11267: dout = 12'h666;
			11268: dout = 12'hfff;
			11269: dout = 12'hddd;
			11270: dout = 12'heee;
			11271: dout = 12'h000;
			11272: dout = 12'h000;
			11273: dout = 12'h000;
			11274: dout = 12'haaa;
			11275: dout = 12'hfff;
			11276: dout = 12'h000;
			11277: dout = 12'hfff;
			11278: dout = 12'h666;
			11279: dout = 12'h000;
			11280: dout = 12'h000;
			11281: dout = 12'h000;
			11282: dout = 12'h000;
			11283: dout = 12'h999;
			11284: dout = 12'hfff;
			11285: dout = 12'hbbb;
			11286: dout = 12'hfff;
			11287: dout = 12'h000;
			11288: dout = 12'h000;
			11289: dout = 12'h000;
			11290: dout = 12'h000;
			11291: dout = 12'h000;
			11292: dout = 12'h000;
			11293: dout = 12'h000;
			11294: dout = 12'h000;
			11295: dout = 12'h000;
			11296: dout = 12'h000;
			11297: dout = 12'h000;
			11298: dout = 12'h000;
			11299: dout = 12'h000;

			11300: dout = 12'h000;
			11301: dout = 12'h000;
			11302: dout = 12'h000;
			11303: dout = 12'h000;
			11304: dout = 12'h000;
			11305: dout = 12'h000;
			11306: dout = 12'h000;
			11307: dout = 12'h000;
			11308: dout = 12'h000;
			11309: dout = 12'h000;
			11310: dout = 12'h000;
			11311: dout = 12'h000;
			11312: dout = 12'h888;
			11313: dout = 12'hfff;
			11314: dout = 12'hfee;
			11315: dout = 12'hfff;
			11316: dout = 12'h000;
			11317: dout = 12'h666;
			11318: dout = 12'hfff;
			11319: dout = 12'h877;
			11320: dout = 12'hfff;
			11321: dout = 12'h222;
			11322: dout = 12'h000;
			11323: dout = 12'h000;
			11324: dout = 12'hddd;
			11325: dout = 12'h777;
			11326: dout = 12'h870;
			11327: dout = 12'hfff;
			11328: dout = 12'h666;
			11329: dout = 12'h000;
			11330: dout = 12'h000;
			11331: dout = 12'h000;
			11332: dout = 12'h999;
			11333: dout = 12'hfff;
			11334: dout = 12'h875;
			11335: dout = 12'h543;
			11336: dout = 12'hfff;
			11337: dout = 12'h000;
			11338: dout = 12'h000;
			11339: dout = 12'h000;
			11340: dout = 12'h000;
			11341: dout = 12'h000;
			11342: dout = 12'h000;
			11343: dout = 12'h000;
			11344: dout = 12'h000;
			11345: dout = 12'h000;
			11346: dout = 12'h000;
			11347: dout = 12'h000;
			11348: dout = 12'h000;
			11349: dout = 12'h000;

			11350: dout = 12'h000;
			11351: dout = 12'h000;
			11352: dout = 12'h000;
			11353: dout = 12'h000;
			11354: dout = 12'h000;
			11355: dout = 12'h000;
			11356: dout = 12'h000;
			11357: dout = 12'h000;
			11358: dout = 12'h000;
			11359: dout = 12'h000;
			11360: dout = 12'h000;
			11361: dout = 12'h000;
			11362: dout = 12'h888;
			11363: dout = 12'hfff;
			11364: dout = 12'h110;
			11365: dout = 12'hfff;
			11366: dout = 12'hfff;
			11367: dout = 12'h000;
			11368: dout = 12'hfff;
			11369: dout = 12'h555;
			11370: dout = 12'hdde;
			11371: dout = 12'hfff;
			11372: dout = 12'h111;
			11373: dout = 12'h222;
			11374: dout = 12'hfff;
			11375: dout = 12'h778;
			11376: dout = 12'h770;
			11377: dout = 12'hfff;
			11378: dout = 12'h555;
			11379: dout = 12'h000;
			11380: dout = 12'h000;
			11381: dout = 12'h999;
			11382: dout = 12'hfff;
			11383: dout = 12'h776;
			11384: dout = 12'h980;
			11385: dout = 12'heef;
			11386: dout = 12'hfff;
			11387: dout = 12'h000;
			11388: dout = 12'h000;
			11389: dout = 12'h000;
			11390: dout = 12'h000;
			11391: dout = 12'h000;
			11392: dout = 12'h000;
			11393: dout = 12'h000;
			11394: dout = 12'h000;
			11395: dout = 12'h000;
			11396: dout = 12'h000;
			11397: dout = 12'h000;
			11398: dout = 12'h000;
			11399: dout = 12'h000;

			11400: dout = 12'h000;
			11401: dout = 12'h000;
			11402: dout = 12'h000;
			11403: dout = 12'h000;
			11404: dout = 12'h000;
			11405: dout = 12'h000;
			11406: dout = 12'h000;
			11407: dout = 12'h000;
			11408: dout = 12'h000;
			11409: dout = 12'h000;
			11410: dout = 12'h000;
			11411: dout = 12'h000;
			11412: dout = 12'h000;
			11413: dout = 12'hfff;
			11414: dout = 12'ha98;
			11415: dout = 12'h760;
			11416: dout = 12'heef;
			11417: dout = 12'hfff;
			11418: dout = 12'hfff;
			11419: dout = 12'hbaa;
			11420: dout = 12'h760;
			11421: dout = 12'hdde;
			11422: dout = 12'hfff;
			11423: dout = 12'hfff;
			11424: dout = 12'hbbd;
			11425: dout = 12'hbb1;
			11426: dout = 12'h761;
			11427: dout = 12'hfff;
			11428: dout = 12'h888;
			11429: dout = 12'h111;
			11430: dout = 12'h888;
			11431: dout = 12'hfff;
			11432: dout = 12'h665;
			11433: dout = 12'hff2;
			11434: dout = 12'h665;
			11435: dout = 12'hfff;
			11436: dout = 12'h555;
			11437: dout = 12'h000;
			11438: dout = 12'h000;
			11439: dout = 12'h000;
			11440: dout = 12'h000;
			11441: dout = 12'h000;
			11442: dout = 12'h000;
			11443: dout = 12'h000;
			11444: dout = 12'h000;
			11445: dout = 12'h000;
			11446: dout = 12'h000;
			11447: dout = 12'h000;
			11448: dout = 12'h000;
			11449: dout = 12'h000;

			11450: dout = 12'h000;
			11451: dout = 12'h000;
			11452: dout = 12'h000;
			11453: dout = 12'h000;
			11454: dout = 12'h000;
			11455: dout = 12'h000;
			11456: dout = 12'h000;
			11457: dout = 12'h000;
			11458: dout = 12'h000;
			11459: dout = 12'h000;
			11460: dout = 12'h000;
			11461: dout = 12'h000;
			11462: dout = 12'h000;
			11463: dout = 12'h777;
			11464: dout = 12'hfff;
			11465: dout = 12'h663;
			11466: dout = 12'h992;
			11467: dout = 12'heef;
			11468: dout = 12'hfff;
			11469: dout = 12'hfff;
			11470: dout = 12'h981;
			11471: dout = 12'haa2;
			11472: dout = 12'h779;
			11473: dout = 12'h779;
			11474: dout = 12'hba1;
			11475: dout = 12'hff4;
			11476: dout = 12'hba2;
			11477: dout = 12'hbbd;
			11478: dout = 12'hfff;
			11479: dout = 12'hfff;
			11480: dout = 12'hfff;
			11481: dout = 12'h665;
			11482: dout = 12'hff3;
			11483: dout = 12'h991;
			11484: dout = 12'heef;
			11485: dout = 12'hfff;
			11486: dout = 12'h000;
			11487: dout = 12'h000;
			11488: dout = 12'h000;
			11489: dout = 12'h000;
			11490: dout = 12'h000;
			11491: dout = 12'h000;
			11492: dout = 12'h000;
			11493: dout = 12'h000;
			11494: dout = 12'h000;
			11495: dout = 12'h000;
			11496: dout = 12'h000;
			11497: dout = 12'h000;
			11498: dout = 12'h000;
			11499: dout = 12'h000;

			11500: dout = 12'h000;
			11501: dout = 12'h000;
			11502: dout = 12'h000;
			11503: dout = 12'h000;
			11504: dout = 12'h000;
			11505: dout = 12'h000;
			11506: dout = 12'h000;
			11507: dout = 12'h000;
			11508: dout = 12'h000;
			11509: dout = 12'h000;
			11510: dout = 12'h000;
			11511: dout = 12'h000;
			11512: dout = 12'h000;
			11513: dout = 12'h000;
			11514: dout = 12'heee;
			11515: dout = 12'hdcd;
			11516: dout = 12'hbb1;
			11517: dout = 12'h981;
			11518: dout = 12'h776;
			11519: dout = 12'h778;
			11520: dout = 12'hcb2;
			11521: dout = 12'hff4;
			11522: dout = 12'hfe3;
			11523: dout = 12'hfe3;
			11524: dout = 12'hff4;
			11525: dout = 12'hfe4;
			11526: dout = 12'hff4;
			11527: dout = 12'hba2;
			11528: dout = 12'h651;
			11529: dout = 12'h661;
			11530: dout = 12'h551;
			11531: dout = 12'hfe3;
			11532: dout = 12'hff4;
			11533: dout = 12'h766;
			11534: dout = 12'hfff;
			11535: dout = 12'h444;
			11536: dout = 12'h000;
			11537: dout = 12'h000;
			11538: dout = 12'h000;
			11539: dout = 12'h000;
			11540: dout = 12'h000;
			11541: dout = 12'h000;
			11542: dout = 12'h000;
			11543: dout = 12'h000;
			11544: dout = 12'h000;
			11545: dout = 12'h000;
			11546: dout = 12'h000;
			11547: dout = 12'h000;
			11548: dout = 12'h000;
			11549: dout = 12'h000;

			11550: dout = 12'h000;
			11551: dout = 12'h000;
			11552: dout = 12'h000;
			11553: dout = 12'h000;
			11554: dout = 12'h000;
			11555: dout = 12'h000;
			11556: dout = 12'h000;
			11557: dout = 12'h000;
			11558: dout = 12'h000;
			11559: dout = 12'h000;
			11560: dout = 12'h555;
			11561: dout = 12'hddd;
			11562: dout = 12'hccc;
			11563: dout = 12'hbcc;
			11564: dout = 12'hccd;
			11565: dout = 12'hfff;
			11566: dout = 12'h665;
			11567: dout = 12'hff4;
			11568: dout = 12'hfe3;
			11569: dout = 12'hee3;
			11570: dout = 12'hff4;
			11571: dout = 12'hfe4;
			11572: dout = 12'hfe4;
			11573: dout = 12'hff4;
			11574: dout = 12'hff4;
			11575: dout = 12'hff4;
			11576: dout = 12'hff4;
			11577: dout = 12'hff4;
			11578: dout = 12'hff4;
			11579: dout = 12'hff4;
			11580: dout = 12'hff4;
			11581: dout = 12'hfe4;
			11582: dout = 12'hff4;
			11583: dout = 12'h766;
			11584: dout = 12'hfff;
			11585: dout = 12'h000;
			11586: dout = 12'h000;
			11587: dout = 12'h000;
			11588: dout = 12'h000;
			11589: dout = 12'h000;
			11590: dout = 12'h000;
			11591: dout = 12'h000;
			11592: dout = 12'h000;
			11593: dout = 12'h000;
			11594: dout = 12'h000;
			11595: dout = 12'h000;
			11596: dout = 12'h000;
			11597: dout = 12'h000;
			11598: dout = 12'h000;
			11599: dout = 12'h000;

			11600: dout = 12'h000;
			11601: dout = 12'h000;
			11602: dout = 12'h000;
			11603: dout = 12'h000;
			11604: dout = 12'h000;
			11605: dout = 12'h000;
			11606: dout = 12'h000;
			11607: dout = 12'h000;
			11608: dout = 12'h555;
			11609: dout = 12'hbbb;
			11610: dout = 12'hfff;
			11611: dout = 12'hbbb;
			11612: dout = 12'haaa;
			11613: dout = 12'haaa;
			11614: dout = 12'hfff;
			11615: dout = 12'hfff;
			11616: dout = 12'h665;
			11617: dout = 12'hff4;
			11618: dout = 12'hff4;
			11619: dout = 12'hff4;
			11620: dout = 12'hfe4;
			11621: dout = 12'hfe4;
			11622: dout = 12'hff4;
			11623: dout = 12'h753;
			11624: dout = 12'h644;
			11625: dout = 12'h744;
			11626: dout = 12'h212;
			11627: dout = 12'hcc3;
			11628: dout = 12'hff4;
			11629: dout = 12'hfe4;
			11630: dout = 12'hfe4;
			11631: dout = 12'hfe4;
			11632: dout = 12'hff4;
			11633: dout = 12'h666;
			11634: dout = 12'hfff;
			11635: dout = 12'h333;
			11636: dout = 12'h000;
			11637: dout = 12'h000;
			11638: dout = 12'h000;
			11639: dout = 12'h000;
			11640: dout = 12'h000;
			11641: dout = 12'h000;
			11642: dout = 12'h000;
			11643: dout = 12'h000;
			11644: dout = 12'h000;
			11645: dout = 12'h000;
			11646: dout = 12'h000;
			11647: dout = 12'h000;
			11648: dout = 12'h000;
			11649: dout = 12'h000;

			11650: dout = 12'h000;
			11651: dout = 12'h000;
			11652: dout = 12'h000;
			11653: dout = 12'h000;
			11654: dout = 12'h000;
			11655: dout = 12'h000;
			11656: dout = 12'h000;
			11657: dout = 12'heee;
			11658: dout = 12'hfff;
			11659: dout = 12'hbbb;
			11660: dout = 12'h677;
			11661: dout = 12'h421;
			11662: dout = 12'h533;
			11663: dout = 12'h532;
			11664: dout = 12'h644;
			11665: dout = 12'hfff;
			11666: dout = 12'h775;
			11667: dout = 12'hbb2;
			11668: dout = 12'h634;
			11669: dout = 12'h644;
			11670: dout = 12'hdd3;
			11671: dout = 12'hff4;
			11672: dout = 12'h753;
			11673: dout = 12'he66;
			11674: dout = 12'he65;
			11675: dout = 12'he65;
			11676: dout = 12'he66;
			11677: dout = 12'h945;
			11678: dout = 12'hcc3;
			11679: dout = 12'hff4;
			11680: dout = 12'hff4;
			11681: dout = 12'hff4;
			11682: dout = 12'hff4;
			11683: dout = 12'hcb2;
			11684: dout = 12'hbbb;
			11685: dout = 12'hfff;
			11686: dout = 12'h333;
			11687: dout = 12'h000;
			11688: dout = 12'h222;
			11689: dout = 12'hbbb;
			11690: dout = 12'h999;
			11691: dout = 12'h000;
			11692: dout = 12'h000;
			11693: dout = 12'h000;
			11694: dout = 12'h000;
			11695: dout = 12'h000;
			11696: dout = 12'h000;
			11697: dout = 12'h000;
			11698: dout = 12'h000;
			11699: dout = 12'h000;

			11700: dout = 12'h000;
			11701: dout = 12'h000;
			11702: dout = 12'h000;
			11703: dout = 12'h000;
			11704: dout = 12'h000;
			11705: dout = 12'h000;
			11706: dout = 12'h000;
			11707: dout = 12'hfff;
			11708: dout = 12'h222;
			11709: dout = 12'h733;
			11710: dout = 12'hd76;
			11711: dout = 12'he66;
			11712: dout = 12'hf66;
			11713: dout = 12'he66;
			11714: dout = 12'he65;
			11715: dout = 12'h744;
			11716: dout = 12'h661;
			11717: dout = 12'hb56;
			11718: dout = 12'he66;
			11719: dout = 12'he66;
			11720: dout = 12'h855;
			11721: dout = 12'h432;
			11722: dout = 12'he66;
			11723: dout = 12'hd32;
			11724: dout = 12'he32;
			11725: dout = 12'he32;
			11726: dout = 12'hd32;
			11727: dout = 12'hf65;
			11728: dout = 12'h000;
			11729: dout = 12'h744;
			11730: dout = 12'h644;
			11731: dout = 12'h644;
			11732: dout = 12'h872;
			11733: dout = 12'hcc3;
			11734: dout = 12'h550;
			11735: dout = 12'heef;
			11736: dout = 12'hfff;
			11737: dout = 12'hddd;
			11738: dout = 12'hfff;
			11739: dout = 12'hccc;
			11740: dout = 12'hfff;
			11741: dout = 12'hfff;
			11742: dout = 12'h999;
			11743: dout = 12'h000;
			11744: dout = 12'h000;
			11745: dout = 12'h000;
			11746: dout = 12'h000;
			11747: dout = 12'h000;
			11748: dout = 12'h000;
			11749: dout = 12'h000;

			11750: dout = 12'h000;
			11751: dout = 12'h000;
			11752: dout = 12'h000;
			11753: dout = 12'h000;
			11754: dout = 12'h000;
			11755: dout = 12'h000;
			11756: dout = 12'h000;
			11757: dout = 12'hfff;
			11758: dout = 12'h111;
			11759: dout = 12'hd54;
			11760: dout = 12'hd43;
			11761: dout = 12'he32;
			11762: dout = 12'ha22;
			11763: dout = 12'hd32;
			11764: dout = 12'he32;
			11765: dout = 12'ha33;
			11766: dout = 12'h855;
			11767: dout = 12'he44;
			11768: dout = 12'hf32;
			11769: dout = 12'he32;
			11770: dout = 12'he54;
			11771: dout = 12'he65;
			11772: dout = 12'he32;
			11773: dout = 12'hf32;
			11774: dout = 12'h511;
			11775: dout = 12'hd32;
			11776: dout = 12'he32;
			11777: dout = 12'he32;
			11778: dout = 12'h533;
			11779: dout = 12'hf66;
			11780: dout = 12'he55;
			11781: dout = 12'hf66;
			11782: dout = 12'h111;
			11783: dout = 12'h734;
			11784: dout = 12'hd77;
			11785: dout = 12'h744;
			11786: dout = 12'h755;
			11787: dout = 12'hfff;
			11788: dout = 12'haaa;
			11789: dout = 12'h311;
			11790: dout = 12'h432;
			11791: dout = 12'h787;
			11792: dout = 12'hfff;
			11793: dout = 12'hfff;
			11794: dout = 12'hfff;
			11795: dout = 12'h888;
			11796: dout = 12'h000;
			11797: dout = 12'h000;
			11798: dout = 12'h000;
			11799: dout = 12'h000;

			11800: dout = 12'h000;
			11801: dout = 12'h000;
			11802: dout = 12'h000;
			11803: dout = 12'h000;
			11804: dout = 12'h000;
			11805: dout = 12'h000;
			11806: dout = 12'h000;
			11807: dout = 12'hfff;
			11808: dout = 12'h121;
			11809: dout = 12'hd32;
			11810: dout = 12'he32;
			11811: dout = 12'hb32;
			11812: dout = 12'h011;
			11813: dout = 12'hb32;
			11814: dout = 12'he32;
			11815: dout = 12'he32;
			11816: dout = 12'hd32;
			11817: dout = 12'hf32;
			11818: dout = 12'h411;
			11819: dout = 12'ha22;
			11820: dout = 12'he32;
			11821: dout = 12'he32;
			11822: dout = 12'hf32;
			11823: dout = 12'h511;
			11824: dout = 12'h231;
			11825: dout = 12'h521;
			11826: dout = 12'hf32;
			11827: dout = 12'he32;
			11828: dout = 12'hd32;
			11829: dout = 12'he32;
			11830: dout = 12'he32;
			11831: dout = 12'hc32;
			11832: dout = 12'h733;
			11833: dout = 12'hf55;
			11834: dout = 12'he32;
			11835: dout = 12'hf54;
			11836: dout = 12'h944;
			11837: dout = 12'h677;
			11838: dout = 12'h532;
			11839: dout = 12'hf66;
			11840: dout = 12'he66;
			11841: dout = 12'hb55;
			11842: dout = 12'h533;
			11843: dout = 12'h543;
			11844: dout = 12'hccc;
			11845: dout = 12'hfff;
			11846: dout = 12'hbbb;
			11847: dout = 12'h000;
			11848: dout = 12'h000;
			11849: dout = 12'h000;

			11850: dout = 12'h000;
			11851: dout = 12'h000;
			11852: dout = 12'h000;
			11853: dout = 12'h000;
			11854: dout = 12'h000;
			11855: dout = 12'h000;
			11856: dout = 12'h000;
			11857: dout = 12'hfff;
			11858: dout = 12'h121;
			11859: dout = 12'hd32;
			11860: dout = 12'he32;
			11861: dout = 12'hb32;
			11862: dout = 12'h521;
			11863: dout = 12'he32;
			11864: dout = 12'hf32;
			11865: dout = 12'h821;
			11866: dout = 12'hf32;
			11867: dout = 12'h721;
			11868: dout = 12'h121;
			11869: dout = 12'h922;
			11870: dout = 12'he32;
			11871: dout = 12'he32;
			11872: dout = 12'hc32;
			11873: dout = 12'h121;
			11874: dout = 12'hff4;
			11875: dout = 12'h000;
			11876: dout = 12'hf32;
			11877: dout = 12'he32;
			11878: dout = 12'he32;
			11879: dout = 12'he32;
			11880: dout = 12'he32;
			11881: dout = 12'hd32;
			11882: dout = 12'he32;
			11883: dout = 12'he32;
			11884: dout = 12'he32;
			11885: dout = 12'he32;
			11886: dout = 12'h111;
			11887: dout = 12'h410;
			11888: dout = 12'hf43;
			11889: dout = 12'he32;
			11890: dout = 12'hd32;
			11891: dout = 12'he44;
			11892: dout = 12'hf76;
			11893: dout = 12'h421;
			11894: dout = 12'h000;
			11895: dout = 12'hfff;
			11896: dout = 12'hbbb;
			11897: dout = 12'h000;
			11898: dout = 12'h000;
			11899: dout = 12'h000;

			11900: dout = 12'h000;
			11901: dout = 12'h000;
			11902: dout = 12'h000;
			11903: dout = 12'h000;
			11904: dout = 12'h000;
			11905: dout = 12'h000;
			11906: dout = 12'h000;
			11907: dout = 12'hfff;
			11908: dout = 12'h111;
			11909: dout = 12'h621;
			11910: dout = 12'he32;
			11911: dout = 12'he32;
			11912: dout = 12'he32;
			11913: dout = 12'he32;
			11914: dout = 12'h932;
			11915: dout = 12'h311;
			11916: dout = 12'hf32;
			11917: dout = 12'h742;
			11918: dout = 12'h672;
			11919: dout = 12'h922;
			11920: dout = 12'he32;
			11921: dout = 12'hf32;
			11922: dout = 12'h511;
			11923: dout = 12'haa3;
			11924: dout = 12'hef4;
			11925: dout = 12'h711;
			11926: dout = 12'he32;
			11927: dout = 12'he32;
			11928: dout = 12'he32;
			11929: dout = 12'hc32;
			11930: dout = 12'he32;
			11931: dout = 12'he32;
			11932: dout = 12'hc32;
			11933: dout = 12'he32;
			11934: dout = 12'hf32;
			11935: dout = 12'h821;
			11936: dout = 12'h521;
			11937: dout = 12'hf32;
			11938: dout = 12'he32;
			11939: dout = 12'he32;
			11940: dout = 12'he32;
			11941: dout = 12'hd32;
			11942: dout = 12'h410;
			11943: dout = 12'h222;
			11944: dout = 12'hbba;
			11945: dout = 12'hfff;
			11946: dout = 12'h000;
			11947: dout = 12'h000;
			11948: dout = 12'h000;
			11949: dout = 12'h000;

			11950: dout = 12'h000;
			11951: dout = 12'h000;
			11952: dout = 12'h000;
			11953: dout = 12'h000;
			11954: dout = 12'h000;
			11955: dout = 12'h000;
			11956: dout = 12'h000;
			11957: dout = 12'hfff;
			11958: dout = 12'h999;
			11959: dout = 12'h510;
			11960: dout = 12'hf32;
			11961: dout = 12'he32;
			11962: dout = 12'he32;
			11963: dout = 12'hf32;
			11964: dout = 12'hc32;
			11965: dout = 12'h721;
			11966: dout = 12'hf32;
			11967: dout = 12'h631;
			11968: dout = 12'h552;
			11969: dout = 12'ha22;
			11970: dout = 12'hf32;
			11971: dout = 12'he32;
			11972: dout = 12'h711;
			11973: dout = 12'h672;
			11974: dout = 12'h621;
			11975: dout = 12'hf32;
			11976: dout = 12'he32;
			11977: dout = 12'he32;
			11978: dout = 12'hd32;
			11979: dout = 12'h621;
			11980: dout = 12'hf32;
			11981: dout = 12'he32;
			11982: dout = 12'h521;
			11983: dout = 12'hf32;
			11984: dout = 12'hb32;
			11985: dout = 12'h011;
			11986: dout = 12'hd32;
			11987: dout = 12'he32;
			11988: dout = 12'he32;
			11989: dout = 12'hf32;
			11990: dout = 12'hb21;
			11991: dout = 12'h000;
			11992: dout = 12'haaa;
			11993: dout = 12'hfff;
			11994: dout = 12'hfff;
			11995: dout = 12'h666;
			11996: dout = 12'h000;
			11997: dout = 12'h000;
			11998: dout = 12'h000;
			11999: dout = 12'h000;

			12000: dout = 12'h000;
			12001: dout = 12'h000;
			12002: dout = 12'h000;
			12003: dout = 12'h000;
			12004: dout = 12'h000;
			12005: dout = 12'h000;
			12006: dout = 12'h000;
			12007: dout = 12'hbbb;
			12008: dout = 12'hbbb;
			12009: dout = 12'h000;
			12010: dout = 12'hd32;
			12011: dout = 12'he32;
			12012: dout = 12'hc32;
			12013: dout = 12'h211;
			12014: dout = 12'hc32;
			12015: dout = 12'hf32;
			12016: dout = 12'he32;
			12017: dout = 12'hb22;
			12018: dout = 12'h411;
			12019: dout = 12'hf32;
			12020: dout = 12'ha22;
			12021: dout = 12'he32;
			12022: dout = 12'he32;
			12023: dout = 12'ha21;
			12024: dout = 12'hd32;
			12025: dout = 12'hd32;
			12026: dout = 12'ha22;
			12027: dout = 12'hf32;
			12028: dout = 12'h621;
			12029: dout = 12'h621;
			12030: dout = 12'hf42;
			12031: dout = 12'h211;
			12032: dout = 12'hb32;
			12033: dout = 12'hf32;
			12034: dout = 12'hb32;
			12035: dout = 12'hb32;
			12036: dout = 12'hf32;
			12037: dout = 12'he32;
			12038: dout = 12'hf32;
			12039: dout = 12'ha21;
			12040: dout = 12'h344;
			12041: dout = 12'heee;
			12042: dout = 12'hfff;
			12043: dout = 12'haaa;
			12044: dout = 12'h000;
			12045: dout = 12'h000;
			12046: dout = 12'h000;
			12047: dout = 12'h000;
			12048: dout = 12'h000;
			12049: dout = 12'h000;

			12050: dout = 12'h000;
			12051: dout = 12'h000;
			12052: dout = 12'h000;
			12053: dout = 12'h000;
			12054: dout = 12'h000;
			12055: dout = 12'h000;
			12056: dout = 12'h000;
			12057: dout = 12'haaa;
			12058: dout = 12'hfff;
			12059: dout = 12'h111;
			12060: dout = 12'hd32;
			12061: dout = 12'he32;
			12062: dout = 12'hb32;
			12063: dout = 12'h011;
			12064: dout = 12'hc32;
			12065: dout = 12'he32;
			12066: dout = 12'he32;
			12067: dout = 12'he32;
			12068: dout = 12'hf42;
			12069: dout = 12'h621;
			12070: dout = 12'h311;
			12071: dout = 12'hf42;
			12072: dout = 12'he32;
			12073: dout = 12'hf32;
			12074: dout = 12'he32;
			12075: dout = 12'h111;
			12076: dout = 12'hd32;
			12077: dout = 12'hd32;
			12078: dout = 12'h011;
			12079: dout = 12'h621;
			12080: dout = 12'ha32;
			12081: dout = 12'h421;
			12082: dout = 12'hd32;
			12083: dout = 12'hc32;
			12084: dout = 12'h421;
			12085: dout = 12'hb32;
			12086: dout = 12'hc32;
			12087: dout = 12'hc32;
			12088: dout = 12'ha21;
			12089: dout = 12'h343;
			12090: dout = 12'hfff;
			12091: dout = 12'hfff;
			12092: dout = 12'h777;
			12093: dout = 12'h000;
			12094: dout = 12'h000;
			12095: dout = 12'h000;
			12096: dout = 12'h000;
			12097: dout = 12'h000;
			12098: dout = 12'h000;
			12099: dout = 12'h000;

			12100: dout = 12'h000;
			12101: dout = 12'h000;
			12102: dout = 12'h000;
			12103: dout = 12'h000;
			12104: dout = 12'h000;
			12105: dout = 12'h000;
			12106: dout = 12'h000;
			12107: dout = 12'h111;
			12108: dout = 12'hfff;
			12109: dout = 12'h222;
			12110: dout = 12'h721;
			12111: dout = 12'hf32;
			12112: dout = 12'hb32;
			12113: dout = 12'h922;
			12114: dout = 12'hf32;
			12115: dout = 12'hb32;
			12116: dout = 12'h411;
			12117: dout = 12'he32;
			12118: dout = 12'h621;
			12119: dout = 12'h111;
			12120: dout = 12'h001;
			12121: dout = 12'ha32;
			12122: dout = 12'hd32;
			12123: dout = 12'hd32;
			12124: dout = 12'h211;
			12125: dout = 12'h001;
			12126: dout = 12'h001;
			12127: dout = 12'h001;
			12128: dout = 12'h101;
			12129: dout = 12'h001;
			12130: dout = 12'h001;
			12131: dout = 12'h111;
			12132: dout = 12'h011;
			12133: dout = 12'h921;
			12134: dout = 12'hb32;
			12135: dout = 12'h821;
			12136: dout = 12'h111;
			12137: dout = 12'h000;
			12138: dout = 12'h333;
			12139: dout = 12'hfff;
			12140: dout = 12'heee;
			12141: dout = 12'h000;
			12142: dout = 12'h000;
			12143: dout = 12'h000;
			12144: dout = 12'h000;
			12145: dout = 12'h000;
			12146: dout = 12'h000;
			12147: dout = 12'h000;
			12148: dout = 12'h000;
			12149: dout = 12'h000;

			12150: dout = 12'h000;
			12151: dout = 12'h000;
			12152: dout = 12'h000;
			12153: dout = 12'h000;
			12154: dout = 12'h000;
			12155: dout = 12'h000;
			12156: dout = 12'h000;
			12157: dout = 12'h111;
			12158: dout = 12'hfff;
			12159: dout = 12'h333;
			12160: dout = 12'h411;
			12161: dout = 12'hf32;
			12162: dout = 12'he32;
			12163: dout = 12'he32;
			12164: dout = 12'he32;
			12165: dout = 12'hb22;
			12166: dout = 12'h001;
			12167: dout = 12'h000;
			12168: dout = 12'h221;
			12169: dout = 12'hff4;
			12170: dout = 12'h552;
			12171: dout = 12'h001;
			12172: dout = 12'h011;
			12173: dout = 12'h011;
			12174: dout = 12'h111;
			12175: dout = 12'hcb3;
			12176: dout = 12'hba3;
			12177: dout = 12'hbb3;
			12178: dout = 12'hbb3;
			12179: dout = 12'hba3;
			12180: dout = 12'hbb3;
			12181: dout = 12'h772;
			12182: dout = 12'hb22;
			12183: dout = 12'hf32;
			12184: dout = 12'he32;
			12185: dout = 12'hf32;
			12186: dout = 12'hf32;
			12187: dout = 12'h533;
			12188: dout = 12'hfff;
			12189: dout = 12'hfff;
			12190: dout = 12'h000;
			12191: dout = 12'h000;
			12192: dout = 12'h000;
			12193: dout = 12'h000;
			12194: dout = 12'h000;
			12195: dout = 12'h000;
			12196: dout = 12'h000;
			12197: dout = 12'h000;
			12198: dout = 12'h000;
			12199: dout = 12'h000;

			12200: dout = 12'h000;
			12201: dout = 12'h000;
			12202: dout = 12'h000;
			12203: dout = 12'h000;
			12204: dout = 12'h000;
			12205: dout = 12'h000;
			12206: dout = 12'h000;
			12207: dout = 12'h000;
			12208: dout = 12'hfff;
			12209: dout = 12'hccc;
			12210: dout = 12'h300;
			12211: dout = 12'hf32;
			12212: dout = 12'he32;
			12213: dout = 12'he32;
			12214: dout = 12'hf32;
			12215: dout = 12'h531;
			12216: dout = 12'hcb2;
			12217: dout = 12'h972;
			12218: dout = 12'haa2;
			12219: dout = 12'hff4;
			12220: dout = 12'hff4;
			12221: dout = 12'h552;
			12222: dout = 12'h211;
			12223: dout = 12'h211;
			12224: dout = 12'hee4;
			12225: dout = 12'hff4;
			12226: dout = 12'hff4;
			12227: dout = 12'hff4;
			12228: dout = 12'hff4;
			12229: dout = 12'hff4;
			12230: dout = 12'hff4;
			12231: dout = 12'haa3;
			12232: dout = 12'h101;
			12233: dout = 12'hd32;
			12234: dout = 12'hd32;
			12235: dout = 12'hd32;
			12236: dout = 12'hb21;
			12237: dout = 12'h555;
			12238: dout = 12'hfff;
			12239: dout = 12'h000;
			12240: dout = 12'h000;
			12241: dout = 12'h000;
			12242: dout = 12'h000;
			12243: dout = 12'h000;
			12244: dout = 12'h000;
			12245: dout = 12'h000;
			12246: dout = 12'h000;
			12247: dout = 12'h000;
			12248: dout = 12'h000;
			12249: dout = 12'h000;

			12250: dout = 12'h000;
			12251: dout = 12'h000;
			12252: dout = 12'h000;
			12253: dout = 12'h000;
			12254: dout = 12'h000;
			12255: dout = 12'h000;
			12256: dout = 12'h000;
			12257: dout = 12'h000;
			12258: dout = 12'hbbb;
			12259: dout = 12'hccc;
			12260: dout = 12'h000;
			12261: dout = 12'hc32;
			12262: dout = 12'hf32;
			12263: dout = 12'hc32;
			12264: dout = 12'h311;
			12265: dout = 12'h431;
			12266: dout = 12'ha93;
			12267: dout = 12'hfff;
			12268: dout = 12'hbbc;
			12269: dout = 12'hba2;
			12270: dout = 12'hff4;
			12271: dout = 12'hff4;
			12272: dout = 12'hff4;
			12273: dout = 12'hff4;
			12274: dout = 12'hff4;
			12275: dout = 12'hfe4;
			12276: dout = 12'hfe4;
			12277: dout = 12'hed3;
			12278: dout = 12'hdd3;
			12279: dout = 12'hdc2;
			12280: dout = 12'hff4;
			12281: dout = 12'haa3;
			12282: dout = 12'h001;
			12283: dout = 12'h010;
			12284: dout = 12'h011;
			12285: dout = 12'h010;
			12286: dout = 12'h000;
			12287: dout = 12'hfff;
			12288: dout = 12'heee;
			12289: dout = 12'h000;
			12290: dout = 12'h000;
			12291: dout = 12'h000;
			12292: dout = 12'h000;
			12293: dout = 12'h000;
			12294: dout = 12'h000;
			12295: dout = 12'h000;
			12296: dout = 12'h000;
			12297: dout = 12'h000;
			12298: dout = 12'h000;
			12299: dout = 12'h000;

			12300: dout = 12'h000;
			12301: dout = 12'h000;
			12302: dout = 12'h000;
			12303: dout = 12'h000;
			12304: dout = 12'h000;
			12305: dout = 12'h000;
			12306: dout = 12'h000;
			12307: dout = 12'h000;
			12308: dout = 12'h444;
			12309: dout = 12'hfff;
			12310: dout = 12'h232;
			12311: dout = 12'hc32;
			12312: dout = 12'hd32;
			12313: dout = 12'h111;
			12314: dout = 12'h331;
			12315: dout = 12'h873;
			12316: dout = 12'hfff;
			12317: dout = 12'hfff;
			12318: dout = 12'hfff;
			12319: dout = 12'hbbc;
			12320: dout = 12'hba2;
			12321: dout = 12'hff4;
			12322: dout = 12'hfe3;
			12323: dout = 12'h552;
			12324: dout = 12'haa2;
			12325: dout = 12'hff4;
			12326: dout = 12'hff4;
			12327: dout = 12'h335;
			12328: dout = 12'ha9a;
			12329: dout = 12'h99b;
			12330: dout = 12'h992;
			12331: dout = 12'hff4;
			12332: dout = 12'h772;
			12333: dout = 12'h111;
			12334: dout = 12'h211;
			12335: dout = 12'h100;
			12336: dout = 12'hbbb;
			12337: dout = 12'hfff;
			12338: dout = 12'h444;
			12339: dout = 12'h000;
			12340: dout = 12'h000;
			12341: dout = 12'h000;
			12342: dout = 12'h000;
			12343: dout = 12'h000;
			12344: dout = 12'h000;
			12345: dout = 12'h000;
			12346: dout = 12'h000;
			12347: dout = 12'h000;
			12348: dout = 12'h000;
			12349: dout = 12'h000;

			12350: dout = 12'h000;
			12351: dout = 12'h000;
			12352: dout = 12'h000;
			12353: dout = 12'h000;
			12354: dout = 12'h000;
			12355: dout = 12'h000;
			12356: dout = 12'h000;
			12357: dout = 12'h000;
			12358: dout = 12'h000;
			12359: dout = 12'hfff;
			12360: dout = 12'h322;
			12361: dout = 12'h010;
			12362: dout = 12'h001;
			12363: dout = 12'h330;
			12364: dout = 12'h882;
			12365: dout = 12'hfff;
			12366: dout = 12'hfff;
			12367: dout = 12'h000;
			12368: dout = 12'h777;
			12369: dout = 12'hfff;
			12370: dout = 12'h881;
			12371: dout = 12'hff4;
			12372: dout = 12'h651;
			12373: dout = 12'hfff;
			12374: dout = 12'hccd;
			12375: dout = 12'h991;
			12376: dout = 12'hff3;
			12377: dout = 12'h778;
			12378: dout = 12'hfff;
			12379: dout = 12'hfff;
			12380: dout = 12'hddf;
			12381: dout = 12'h992;
			12382: dout = 12'ha91;
			12383: dout = 12'hfff;
			12384: dout = 12'hfff;
			12385: dout = 12'hfff;
			12386: dout = 12'hfff;
			12387: dout = 12'h555;
			12388: dout = 12'h000;
			12389: dout = 12'h000;
			12390: dout = 12'h000;
			12391: dout = 12'h000;
			12392: dout = 12'h000;
			12393: dout = 12'h000;
			12394: dout = 12'h000;
			12395: dout = 12'h000;
			12396: dout = 12'h000;
			12397: dout = 12'h000;
			12398: dout = 12'h000;
			12399: dout = 12'h000;

			12400: dout = 12'h000;
			12401: dout = 12'h000;
			12402: dout = 12'h000;
			12403: dout = 12'h000;
			12404: dout = 12'h000;
			12405: dout = 12'h000;
			12406: dout = 12'h000;
			12407: dout = 12'h000;
			12408: dout = 12'h000;
			12409: dout = 12'hfff;
			12410: dout = 12'h221;
			12411: dout = 12'h000;
			12412: dout = 12'h320;
			12413: dout = 12'h872;
			12414: dout = 12'hfff;
			12415: dout = 12'hfff;
			12416: dout = 12'h000;
			12417: dout = 12'h000;
			12418: dout = 12'h555;
			12419: dout = 12'hfff;
			12420: dout = 12'h874;
			12421: dout = 12'hfe3;
			12422: dout = 12'h88a;
			12423: dout = 12'hfff;
			12424: dout = 12'hfff;
			12425: dout = 12'hccd;
			12426: dout = 12'hba1;
			12427: dout = 12'h878;
			12428: dout = 12'hfff;
			12429: dout = 12'h000;
			12430: dout = 12'hfff;
			12431: dout = 12'heef;
			12432: dout = 12'h760;
			12433: dout = 12'haa9;
			12434: dout = 12'hfff;
			12435: dout = 12'h333;
			12436: dout = 12'h222;
			12437: dout = 12'h000;
			12438: dout = 12'h000;
			12439: dout = 12'h000;
			12440: dout = 12'h000;
			12441: dout = 12'h000;
			12442: dout = 12'h000;
			12443: dout = 12'h000;
			12444: dout = 12'h000;
			12445: dout = 12'h000;
			12446: dout = 12'h000;
			12447: dout = 12'h000;
			12448: dout = 12'h000;
			12449: dout = 12'h000;

			12450: dout = 12'h000;
			12451: dout = 12'h000;
			12452: dout = 12'h000;
			12453: dout = 12'h000;
			12454: dout = 12'h000;
			12455: dout = 12'h000;
			12456: dout = 12'h000;
			12457: dout = 12'h000;
			12458: dout = 12'h000;
			12459: dout = 12'hfff;
			12460: dout = 12'haaa;
			12461: dout = 12'hcbb;
			12462: dout = 12'hfff;
			12463: dout = 12'hfff;
			12464: dout = 12'hfff;
			12465: dout = 12'h000;
			12466: dout = 12'h000;
			12467: dout = 12'h000;
			12468: dout = 12'h000;
			12469: dout = 12'hfff;
			12470: dout = 12'h766;
			12471: dout = 12'hba2;
			12472: dout = 12'hdde;
			12473: dout = 12'hccc;
			12474: dout = 12'h222;
			12475: dout = 12'hfff;
			12476: dout = 12'h660;
			12477: dout = 12'h878;
			12478: dout = 12'hfff;
			12479: dout = 12'h000;
			12480: dout = 12'h000;
			12481: dout = 12'hfff;
			12482: dout = 12'heee;
			12483: dout = 12'h554;
			12484: dout = 12'hfff;
			12485: dout = 12'h000;
			12486: dout = 12'h000;
			12487: dout = 12'h000;
			12488: dout = 12'h000;
			12489: dout = 12'h000;
			12490: dout = 12'h000;
			12491: dout = 12'h000;
			12492: dout = 12'h000;
			12493: dout = 12'h000;
			12494: dout = 12'h000;
			12495: dout = 12'h000;
			12496: dout = 12'h000;
			12497: dout = 12'h000;
			12498: dout = 12'h000;
			12499: dout = 12'h000;

			12500: dout = 12'h000;
			12501: dout = 12'h000;
			12502: dout = 12'h000;
			12503: dout = 12'h000;
			12504: dout = 12'h000;
			12505: dout = 12'h000;
			12506: dout = 12'h000;
			12507: dout = 12'h000;
			12508: dout = 12'h000;
			12509: dout = 12'h888;
			12510: dout = 12'hfff;
			12511: dout = 12'hfff;
			12512: dout = 12'hddd;
			12513: dout = 12'hccc;
			12514: dout = 12'h000;
			12515: dout = 12'h000;
			12516: dout = 12'h000;
			12517: dout = 12'h000;
			12518: dout = 12'h000;
			12519: dout = 12'hbbb;
			12520: dout = 12'hfff;
			12521: dout = 12'h000;
			12522: dout = 12'hfff;
			12523: dout = 12'h333;
			12524: dout = 12'h000;
			12525: dout = 12'hfff;
			12526: dout = 12'hccd;
			12527: dout = 12'h777;
			12528: dout = 12'hfff;
			12529: dout = 12'h000;
			12530: dout = 12'h000;
			12531: dout = 12'h000;
			12532: dout = 12'hfff;
			12533: dout = 12'hfff;
			12534: dout = 12'heee;
			12535: dout = 12'h000;
			12536: dout = 12'h000;
			12537: dout = 12'h000;
			12538: dout = 12'h000;
			12539: dout = 12'h000;
			12540: dout = 12'h000;
			12541: dout = 12'h000;
			12542: dout = 12'h000;
			12543: dout = 12'h000;
			12544: dout = 12'h000;
			12545: dout = 12'h000;
			12546: dout = 12'h000;
			12547: dout = 12'h000;
			12548: dout = 12'h000;
			12549: dout = 12'h000;

			12550: dout = 12'h000;
			12551: dout = 12'h000;
			12552: dout = 12'h000;
			12553: dout = 12'h000;
			12554: dout = 12'h000;
			12555: dout = 12'h000;
			12556: dout = 12'h000;
			12557: dout = 12'h000;
			12558: dout = 12'h000;
			12559: dout = 12'h000;
			12560: dout = 12'h000;
			12561: dout = 12'h000;
			12562: dout = 12'h000;
			12563: dout = 12'h000;
			12564: dout = 12'h000;
			12565: dout = 12'h000;
			12566: dout = 12'h000;
			12567: dout = 12'h000;
			12568: dout = 12'h000;
			12569: dout = 12'h444;
			12570: dout = 12'hfff;
			12571: dout = 12'ha99;
			12572: dout = 12'hfff;
			12573: dout = 12'h000;
			12574: dout = 12'h000;
			12575: dout = 12'h444;
			12576: dout = 12'hfff;
			12577: dout = 12'h666;
			12578: dout = 12'hfff;
			12579: dout = 12'h000;
			12580: dout = 12'h000;
			12581: dout = 12'h000;
			12582: dout = 12'h000;
			12583: dout = 12'h444;
			12584: dout = 12'h000;
			12585: dout = 12'h000;
			12586: dout = 12'h000;
			12587: dout = 12'h000;
			12588: dout = 12'h000;
			12589: dout = 12'h000;
			12590: dout = 12'h000;
			12591: dout = 12'h000;
			12592: dout = 12'h000;
			12593: dout = 12'h000;
			12594: dout = 12'h000;
			12595: dout = 12'h000;
			12596: dout = 12'h000;
			12597: dout = 12'h000;
			12598: dout = 12'h000;
			12599: dout = 12'h000;

			12600: dout = 12'h000;
			12601: dout = 12'h000;
			12602: dout = 12'h000;
			12603: dout = 12'h000;
			12604: dout = 12'h000;
			12605: dout = 12'h000;
			12606: dout = 12'h000;
			12607: dout = 12'h000;
			12608: dout = 12'h000;
			12609: dout = 12'h000;
			12610: dout = 12'h000;
			12611: dout = 12'h000;
			12612: dout = 12'h000;
			12613: dout = 12'h000;
			12614: dout = 12'h000;
			12615: dout = 12'h000;
			12616: dout = 12'h000;
			12617: dout = 12'h000;
			12618: dout = 12'h000;
			12619: dout = 12'h555;
			12620: dout = 12'hfff;
			12621: dout = 12'h999;
			12622: dout = 12'hddd;
			12623: dout = 12'h000;
			12624: dout = 12'h000;
			12625: dout = 12'h111;
			12626: dout = 12'hfff;
			12627: dout = 12'hfff;
			12628: dout = 12'hccc;
			12629: dout = 12'h000;
			12630: dout = 12'h000;
			12631: dout = 12'h000;
			12632: dout = 12'h000;
			12633: dout = 12'h000;
			12634: dout = 12'h000;
			12635: dout = 12'h000;
			12636: dout = 12'h000;
			12637: dout = 12'h000;
			12638: dout = 12'h000;
			12639: dout = 12'h000;
			12640: dout = 12'h000;
			12641: dout = 12'h000;
			12642: dout = 12'h000;
			12643: dout = 12'h000;
			12644: dout = 12'h000;
			12645: dout = 12'h000;
			12646: dout = 12'h000;
			12647: dout = 12'h000;
			12648: dout = 12'h000;
			12649: dout = 12'h000;

			12650: dout = 12'h000;
			12651: dout = 12'h000;
			12652: dout = 12'h000;
			12653: dout = 12'h000;
			12654: dout = 12'h000;
			12655: dout = 12'h000;
			12656: dout = 12'h000;
			12657: dout = 12'h000;
			12658: dout = 12'h000;
			12659: dout = 12'h000;
			12660: dout = 12'h000;
			12661: dout = 12'h000;
			12662: dout = 12'h000;
			12663: dout = 12'h000;
			12664: dout = 12'h000;
			12665: dout = 12'h000;
			12666: dout = 12'h000;
			12667: dout = 12'h000;
			12668: dout = 12'h000;
			12669: dout = 12'h555;
			12670: dout = 12'hfff;
			12671: dout = 12'h988;
			12672: dout = 12'hddd;
			12673: dout = 12'h000;
			12674: dout = 12'h000;
			12675: dout = 12'h000;
			12676: dout = 12'h111;
			12677: dout = 12'h555;
			12678: dout = 12'h000;
			12679: dout = 12'h000;
			12680: dout = 12'h000;
			12681: dout = 12'h000;
			12682: dout = 12'h000;
			12683: dout = 12'h000;
			12684: dout = 12'h000;
			12685: dout = 12'h000;
			12686: dout = 12'h000;
			12687: dout = 12'h000;
			12688: dout = 12'h000;
			12689: dout = 12'h000;
			12690: dout = 12'h000;
			12691: dout = 12'h000;
			12692: dout = 12'h000;
			12693: dout = 12'h000;
			12694: dout = 12'h000;
			12695: dout = 12'h000;
			12696: dout = 12'h000;
			12697: dout = 12'h000;
			12698: dout = 12'h000;
			12699: dout = 12'h000;

			12700: dout = 12'h000;
			12701: dout = 12'h000;
			12702: dout = 12'h000;
			12703: dout = 12'h000;
			12704: dout = 12'h000;
			12705: dout = 12'h000;
			12706: dout = 12'h000;
			12707: dout = 12'h000;
			12708: dout = 12'h000;
			12709: dout = 12'h000;
			12710: dout = 12'h000;
			12711: dout = 12'h000;
			12712: dout = 12'h000;
			12713: dout = 12'h000;
			12714: dout = 12'h000;
			12715: dout = 12'h000;
			12716: dout = 12'h000;
			12717: dout = 12'h000;
			12718: dout = 12'h000;
			12719: dout = 12'h222;
			12720: dout = 12'hfff;
			12721: dout = 12'hfff;
			12722: dout = 12'haaa;
			12723: dout = 12'h000;
			12724: dout = 12'h000;
			12725: dout = 12'h000;
			12726: dout = 12'h000;
			12727: dout = 12'h000;
			12728: dout = 12'h000;
			12729: dout = 12'h000;
			12730: dout = 12'h000;
			12731: dout = 12'h000;
			12732: dout = 12'h000;
			12733: dout = 12'h000;
			12734: dout = 12'h000;
			12735: dout = 12'h000;
			12736: dout = 12'h000;
			12737: dout = 12'h000;
			12738: dout = 12'h000;
			12739: dout = 12'h000;
			12740: dout = 12'h000;
			12741: dout = 12'h000;
			12742: dout = 12'h000;
			12743: dout = 12'h000;
			12744: dout = 12'h000;
			12745: dout = 12'h000;
			12746: dout = 12'h000;
			12747: dout = 12'h000;
			12748: dout = 12'h000;
			12749: dout = 12'h000;

			12750: dout = 12'h000;
			12751: dout = 12'h000;
			12752: dout = 12'h000;
			12753: dout = 12'h000;
			12754: dout = 12'h000;
			12755: dout = 12'h000;
			12756: dout = 12'h000;
			12757: dout = 12'h000;
			12758: dout = 12'h000;
			12759: dout = 12'h000;
			12760: dout = 12'h000;
			12761: dout = 12'h000;
			12762: dout = 12'h000;
			12763: dout = 12'h000;
			12764: dout = 12'h000;
			12765: dout = 12'h000;
			12766: dout = 12'h000;
			12767: dout = 12'h000;
			12768: dout = 12'h000;
			12769: dout = 12'h000;
			12770: dout = 12'h333;
			12771: dout = 12'h555;
			12772: dout = 12'h000;
			12773: dout = 12'h000;
			12774: dout = 12'h000;
			12775: dout = 12'h000;
			12776: dout = 12'h000;
			12777: dout = 12'h000;
			12778: dout = 12'h000;
			12779: dout = 12'h000;
			12780: dout = 12'h000;
			12781: dout = 12'h000;
			12782: dout = 12'h000;
			12783: dout = 12'h000;
			12784: dout = 12'h000;
			12785: dout = 12'h000;
			12786: dout = 12'h000;
			12787: dout = 12'h000;
			12788: dout = 12'h000;
			12789: dout = 12'h000;
			12790: dout = 12'h000;
			12791: dout = 12'h000;
			12792: dout = 12'h000;
			12793: dout = 12'h000;
			12794: dout = 12'h000;
			12795: dout = 12'h000;
			12796: dout = 12'h000;
			12797: dout = 12'h000;
			12798: dout = 12'h000;
			12799: dout = 12'h000;

			12800: dout = 12'h000;
			12801: dout = 12'h000;
			12802: dout = 12'h000;
			12803: dout = 12'h000;
			12804: dout = 12'h000;
			12805: dout = 12'h000;
			12806: dout = 12'h000;
			12807: dout = 12'h000;
			12808: dout = 12'h000;
			12809: dout = 12'h000;
			12810: dout = 12'h000;
			12811: dout = 12'h000;
			12812: dout = 12'h000;
			12813: dout = 12'h000;
			12814: dout = 12'h000;
			12815: dout = 12'h000;
			12816: dout = 12'h000;
			12817: dout = 12'h000;
			12818: dout = 12'h000;
			12819: dout = 12'h000;
			12820: dout = 12'h000;
			12821: dout = 12'h000;
			12822: dout = 12'h000;
			12823: dout = 12'h000;
			12824: dout = 12'h000;
			12825: dout = 12'h000;
			12826: dout = 12'h000;
			12827: dout = 12'h000;
			12828: dout = 12'h000;
			12829: dout = 12'h000;
			12830: dout = 12'h000;
			12831: dout = 12'h000;
			12832: dout = 12'h000;
			12833: dout = 12'h000;
			12834: dout = 12'h000;
			12835: dout = 12'h000;
			12836: dout = 12'h000;
			12837: dout = 12'h000;
			12838: dout = 12'h000;
			12839: dout = 12'h000;
			12840: dout = 12'h000;
			12841: dout = 12'h000;
			12842: dout = 12'h000;
			12843: dout = 12'h000;
			12844: dout = 12'h000;
			12845: dout = 12'h000;
			12846: dout = 12'h000;
			12847: dout = 12'h000;
			12848: dout = 12'h000;
			12849: dout = 12'h000;

			12850: dout = 12'h000;
			12851: dout = 12'h000;
			12852: dout = 12'h000;
			12853: dout = 12'h000;
			12854: dout = 12'h000;
			12855: dout = 12'h000;
			12856: dout = 12'h000;
			12857: dout = 12'h000;
			12858: dout = 12'h000;
			12859: dout = 12'h000;
			12860: dout = 12'h000;
			12861: dout = 12'h000;
			12862: dout = 12'h000;
			12863: dout = 12'h000;
			12864: dout = 12'h000;
			12865: dout = 12'h000;
			12866: dout = 12'h000;
			12867: dout = 12'h000;
			12868: dout = 12'h000;
			12869: dout = 12'h000;
			12870: dout = 12'h000;
			12871: dout = 12'h000;
			12872: dout = 12'h000;
			12873: dout = 12'h000;
			12874: dout = 12'h000;
			12875: dout = 12'h000;
			12876: dout = 12'h000;
			12877: dout = 12'h000;
			12878: dout = 12'h000;
			12879: dout = 12'h000;
			12880: dout = 12'h000;
			12881: dout = 12'h000;
			12882: dout = 12'h000;
			12883: dout = 12'h000;
			12884: dout = 12'h000;
			12885: dout = 12'h000;
			12886: dout = 12'h000;
			12887: dout = 12'h000;
			12888: dout = 12'h000;
			12889: dout = 12'h000;
			12890: dout = 12'h000;
			12891: dout = 12'h000;
			12892: dout = 12'h000;
			12893: dout = 12'h000;
			12894: dout = 12'h000;
			12895: dout = 12'h000;
			12896: dout = 12'h000;
			12897: dout = 12'h000;
			12898: dout = 12'h000;
			12899: dout = 12'h000;

			12900: dout = 12'h000;
			12901: dout = 12'h000;
			12902: dout = 12'h000;
			12903: dout = 12'h000;
			12904: dout = 12'h000;
			12905: dout = 12'h000;
			12906: dout = 12'h000;
			12907: dout = 12'h000;
			12908: dout = 12'h000;
			12909: dout = 12'h000;
			12910: dout = 12'h000;
			12911: dout = 12'h000;
			12912: dout = 12'h000;
			12913: dout = 12'h000;
			12914: dout = 12'h000;
			12915: dout = 12'h000;
			12916: dout = 12'h000;
			12917: dout = 12'h000;
			12918: dout = 12'h000;
			12919: dout = 12'h000;
			12920: dout = 12'h000;
			12921: dout = 12'h000;
			12922: dout = 12'h000;
			12923: dout = 12'h000;
			12924: dout = 12'h000;
			12925: dout = 12'h000;
			12926: dout = 12'h000;
			12927: dout = 12'h000;
			12928: dout = 12'h000;
			12929: dout = 12'h000;
			12930: dout = 12'h000;
			12931: dout = 12'h000;
			12932: dout = 12'h000;
			12933: dout = 12'h000;
			12934: dout = 12'h000;
			12935: dout = 12'h000;
			12936: dout = 12'h000;
			12937: dout = 12'h000;
			12938: dout = 12'h000;
			12939: dout = 12'h000;
			12940: dout = 12'h000;
			12941: dout = 12'h000;
			12942: dout = 12'h000;
			12943: dout = 12'h000;
			12944: dout = 12'h000;
			12945: dout = 12'h000;
			12946: dout = 12'h000;
			12947: dout = 12'h000;
			12948: dout = 12'h000;
			12949: dout = 12'h000;

			12950: dout = 12'h000;
			12951: dout = 12'h000;
			12952: dout = 12'h000;
			12953: dout = 12'h000;
			12954: dout = 12'h000;
			12955: dout = 12'h000;
			12956: dout = 12'h000;
			12957: dout = 12'h000;
			12958: dout = 12'h000;
			12959: dout = 12'h000;
			12960: dout = 12'h000;
			12961: dout = 12'h000;
			12962: dout = 12'h000;
			12963: dout = 12'h000;
			12964: dout = 12'h000;
			12965: dout = 12'h000;
			12966: dout = 12'h000;
			12967: dout = 12'h000;
			12968: dout = 12'h000;
			12969: dout = 12'h000;
			12970: dout = 12'h000;
			12971: dout = 12'h000;
			12972: dout = 12'h000;
			12973: dout = 12'h000;
			12974: dout = 12'h000;
			12975: dout = 12'h000;
			12976: dout = 12'h000;
			12977: dout = 12'h000;
			12978: dout = 12'h000;
			12979: dout = 12'h000;
			12980: dout = 12'h000;
			12981: dout = 12'h000;
			12982: dout = 12'h000;
			12983: dout = 12'h000;
			12984: dout = 12'h000;
			12985: dout = 12'h000;
			12986: dout = 12'h000;
			12987: dout = 12'h000;
			12988: dout = 12'h000;
			12989: dout = 12'h000;
			12990: dout = 12'h000;
			12991: dout = 12'h000;
			12992: dout = 12'h000;
			12993: dout = 12'h000;
			12994: dout = 12'h000;
			12995: dout = 12'h000;
			12996: dout = 12'h000;
			12997: dout = 12'h000;
			12998: dout = 12'h000;
			12999: dout = 12'h000;

			13000: dout = 12'h000;
			13001: dout = 12'h000;
			13002: dout = 12'h000;
			13003: dout = 12'h000;
			13004: dout = 12'h000;
			13005: dout = 12'h000;
			13006: dout = 12'h000;
			13007: dout = 12'h000;
			13008: dout = 12'h000;
			13009: dout = 12'h000;
			13010: dout = 12'h000;
			13011: dout = 12'h000;
			13012: dout = 12'h000;
			13013: dout = 12'h000;
			13014: dout = 12'h000;
			13015: dout = 12'h000;
			13016: dout = 12'h000;
			13017: dout = 12'h000;
			13018: dout = 12'h000;
			13019: dout = 12'h000;
			13020: dout = 12'h000;
			13021: dout = 12'h000;
			13022: dout = 12'h000;
			13023: dout = 12'h000;
			13024: dout = 12'h000;
			13025: dout = 12'h000;
			13026: dout = 12'h000;
			13027: dout = 12'h000;
			13028: dout = 12'h000;
			13029: dout = 12'h000;
			13030: dout = 12'h000;
			13031: dout = 12'h000;
			13032: dout = 12'h000;
			13033: dout = 12'h000;
			13034: dout = 12'h000;
			13035: dout = 12'h000;
			13036: dout = 12'h000;
			13037: dout = 12'h000;
			13038: dout = 12'h000;
			13039: dout = 12'h000;
			13040: dout = 12'h000;
			13041: dout = 12'h000;
			13042: dout = 12'h000;
			13043: dout = 12'h000;
			13044: dout = 12'h000;
			13045: dout = 12'h000;
			13046: dout = 12'h000;
			13047: dout = 12'h000;
			13048: dout = 12'h000;
			13049: dout = 12'h000;

			13050: dout = 12'h000;
			13051: dout = 12'h000;
			13052: dout = 12'h000;
			13053: dout = 12'h000;
			13054: dout = 12'h000;
			13055: dout = 12'h000;
			13056: dout = 12'h000;
			13057: dout = 12'h000;
			13058: dout = 12'h000;
			13059: dout = 12'h000;
			13060: dout = 12'h000;
			13061: dout = 12'h000;
			13062: dout = 12'h000;
			13063: dout = 12'h000;
			13064: dout = 12'h000;
			13065: dout = 12'h000;
			13066: dout = 12'h000;
			13067: dout = 12'h000;
			13068: dout = 12'h000;
			13069: dout = 12'h000;
			13070: dout = 12'h000;
			13071: dout = 12'h000;
			13072: dout = 12'h000;
			13073: dout = 12'h000;
			13074: dout = 12'h000;
			13075: dout = 12'h000;
			13076: dout = 12'h000;
			13077: dout = 12'h000;
			13078: dout = 12'h000;
			13079: dout = 12'h000;
			13080: dout = 12'h000;
			13081: dout = 12'h000;
			13082: dout = 12'h000;
			13083: dout = 12'h000;
			13084: dout = 12'h000;
			13085: dout = 12'h000;
			13086: dout = 12'h000;
			13087: dout = 12'h000;
			13088: dout = 12'h000;
			13089: dout = 12'h000;
			13090: dout = 12'h000;
			13091: dout = 12'h000;
			13092: dout = 12'h000;
			13093: dout = 12'h000;
			13094: dout = 12'h000;
			13095: dout = 12'h000;
			13096: dout = 12'h000;
			13097: dout = 12'h000;
			13098: dout = 12'h000;
			13099: dout = 12'h000;
			13100: dout = 12'h000;
			13101: dout = 12'h000;
			13102: dout = 12'h000;
			13103: dout = 12'h000;
			13104: dout = 12'h000;
			13105: dout = 12'h000;
			13106: dout = 12'h000;
			13107: dout = 12'h000;
			13108: dout = 12'h000;
			13109: dout = 12'h000;
			13110: dout = 12'h000;
			13111: dout = 12'h000;
			13112: dout = 12'h000;
			13113: dout = 12'h000;
			13114: dout = 12'h000;
			13115: dout = 12'h000;
			13116: dout = 12'h000;
			13117: dout = 12'h000;
			13118: dout = 12'h000;
			13119: dout = 12'h000;
			13120: dout = 12'h000;
			13121: dout = 12'h000;
			13122: dout = 12'h000;
			13123: dout = 12'h000;
			13124: dout = 12'h000;
			13125: dout = 12'h000;
			13126: dout = 12'h000;
			13127: dout = 12'h000;
			13128: dout = 12'h000;
			13129: dout = 12'h000;
			13130: dout = 12'h000;
			13131: dout = 12'h000;
			13132: dout = 12'h000;
			13133: dout = 12'h000;
			13134: dout = 12'h000;
			13135: dout = 12'h000;
			13136: dout = 12'h000;
			13137: dout = 12'h000;
			13138: dout = 12'h000;
			13139: dout = 12'h000;
			13140: dout = 12'h000;
			13141: dout = 12'h000;
			13142: dout = 12'h000;
			13143: dout = 12'h000;
			13144: dout = 12'h000;
			13145: dout = 12'h000;
			13146: dout = 12'h000;
			13147: dout = 12'h000;
			13148: dout = 12'h000;
			13149: dout = 12'h000;
			13150: dout = 12'h000;
			13151: dout = 12'h000;
			13152: dout = 12'h000;
			13153: dout = 12'h000;
			13154: dout = 12'h000;
			13155: dout = 12'h000;
			13156: dout = 12'h000;
			13157: dout = 12'h000;
			13158: dout = 12'h000;
			13159: dout = 12'h000;
			13160: dout = 12'h000;
			13161: dout = 12'h000;
			13162: dout = 12'h000;
			13163: dout = 12'h000;
			13164: dout = 12'h000;
			13165: dout = 12'h000;
			13166: dout = 12'h000;
			13167: dout = 12'h000;
			13168: dout = 12'h000;
			13169: dout = 12'h000;
			13170: dout = 12'h000;
			13171: dout = 12'h000;
			13172: dout = 12'h000;
			13173: dout = 12'h000;
			13174: dout = 12'h000;
			13175: dout = 12'h000;
			13176: dout = 12'h000;
			13177: dout = 12'h000;
			13178: dout = 12'h000;
			13179: dout = 12'h000;
			13180: dout = 12'h000;
			13181: dout = 12'h000;
			13182: dout = 12'h000;
			13183: dout = 12'h000;
			13184: dout = 12'h000;
			13185: dout = 12'h000;
			13186: dout = 12'h000;
			13187: dout = 12'h000;
			13188: dout = 12'h000;
			13189: dout = 12'h000;
			13190: dout = 12'h000;
			13191: dout = 12'h000;
			13192: dout = 12'h000;
			13193: dout = 12'h000;
			13194: dout = 12'h000;
			13195: dout = 12'h000;

			13196: dout = 12'h000;
			13197: dout = 12'h000;
			13198: dout = 12'haaa;
			13199: dout = 12'hccc;
			13200: dout = 12'hccc;
			13201: dout = 12'hccc;
			13202: dout = 12'hddd;
			13203: dout = 12'hddd;
			13204: dout = 12'h777;
			13205: dout = 12'h444;
			13206: dout = 12'h222;
			13207: dout = 12'h000;
			13208: dout = 12'h000;
			13209: dout = 12'h000;
			13210: dout = 12'h000;
			13211: dout = 12'h000;
			13212: dout = 12'h000;
			13213: dout = 12'h000;
			13214: dout = 12'h000;
			13215: dout = 12'h000;
			13216: dout = 12'h000;
			13217: dout = 12'h000;
			13218: dout = 12'h000;
			13219: dout = 12'h000;
			13220: dout = 12'h000;
			13221: dout = 12'h000;
			13222: dout = 12'h000;
			13223: dout = 12'h000;
			13224: dout = 12'h000;
			13225: dout = 12'h000;
			13226: dout = 12'h000;
			13227: dout = 12'h888;
			13228: dout = 12'hfff;
			13229: dout = 12'hfff;
			13230: dout = 12'hfff;
			13231: dout = 12'h888;
			13232: dout = 12'h000;
			13233: dout = 12'h000;
			13234: dout = 12'h000;
			13235: dout = 12'h000;
			13236: dout = 12'h000;
			13237: dout = 12'h000;
			13238: dout = 12'h000;
			13239: dout = 12'h000;
			13240: dout = 12'h000;
			13241: dout = 12'h000;
			13242: dout = 12'h000;
			13243: dout = 12'h000;
			13244: dout = 12'h000;
			13245: dout = 12'h000;
			13246: dout = 12'h000;
			13247: dout = 12'h000;
			13248: dout = 12'h000;
			13249: dout = 12'h000;
			13250: dout = 12'h000;
			13251: dout = 12'h000;
			13252: dout = 12'h000;
			13253: dout = 12'h000;
			13254: dout = 12'h445;
			13255: dout = 12'hddd;
			13256: dout = 12'hbbb;
			13257: dout = 12'h555;
			13258: dout = 12'h444;
			13259: dout = 12'h222;
			13260: dout = 12'h000;
			13261: dout = 12'h000;
			13262: dout = 12'h000;
			13263: dout = 12'h000;
			13264: dout = 12'h000;
			13265: dout = 12'h000;
			13266: dout = 12'h000;
			13267: dout = 12'h000;
			13268: dout = 12'h122;
			13269: dout = 12'hccc;
			13270: dout = 12'hccc;
			13271: dout = 12'hccc;
			13272: dout = 12'hccc;
			13273: dout = 12'hddd;
			13274: dout = 12'hddd;
			13275: dout = 12'h444;
			13276: dout = 12'h444;
			13277: dout = 12'h000;
			13278: dout = 12'h000;
			13279: dout = 12'h000;
			13280: dout = 12'h000;
			13281: dout = 12'h000;
			13282: dout = 12'h000;
			13283: dout = 12'h000;
			13284: dout = 12'h000;
			13285: dout = 12'h000;
			13286: dout = 12'h000;
			13287: dout = 12'h000;
			13288: dout = 12'h111;
			13289: dout = 12'h777;
			13290: dout = 12'h555;
			13291: dout = 12'h444;
			13292: dout = 12'h222;
			13293: dout = 12'h000;
			13294: dout = 12'h010;
			13295: dout = 12'h777;
			13296: dout = 12'h555;
			13297: dout = 12'h444;
			13298: dout = 12'h222;
			13299: dout = 12'h000;
			13300: dout = 12'h000;
			13301: dout = 12'h000;
			13302: dout = 12'h000;
			13303: dout = 12'h000;
			13304: dout = 12'h000;
			13305: dout = 12'h000;
			13306: dout = 12'h000;
			13307: dout = 12'h000;
			13308: dout = 12'h000;
			13309: dout = 12'h000;
			13310: dout = 12'h000;
			13311: dout = 12'h000;
			13312: dout = 12'h000;
			13313: dout = 12'h000;
			13314: dout = 12'h000;
			13315: dout = 12'h000;
			13316: dout = 12'h000;
			13317: dout = 12'h000;
			13318: dout = 12'h000;
			13319: dout = 12'h000;
			13320: dout = 12'h000;
			13321: dout = 12'h000;
			13322: dout = 12'h000;
			13323: dout = 12'h000;
			13324: dout = 12'h000;
			13325: dout = 12'h000;
			13326: dout = 12'h000;
			13327: dout = 12'h000;
			13328: dout = 12'h000;
			13329: dout = 12'h000;
			13330: dout = 12'h000;
			13331: dout = 12'h000;
			13332: dout = 12'h000;
			13333: dout = 12'h000;
			13334: dout = 12'h000;
			13335: dout = 12'h000;
			13336: dout = 12'h000;
			13337: dout = 12'h000;
			13338: dout = 12'h000;
			13339: dout = 12'h000;
			13340: dout = 12'h000;
			13341: dout = 12'h000;

			13342: dout = 12'h000;
			13343: dout = 12'hfff;
			13344: dout = 12'hfff;
			13345: dout = 12'haab;
			13346: dout = 12'habb;
			13347: dout = 12'hbcc;
			13348: dout = 12'h9aa;
			13349: dout = 12'h9aa;
			13350: dout = 12'hfff;
			13351: dout = 12'hfff;
			13352: dout = 12'hfff;
			13353: dout = 12'hddd;
			13354: dout = 12'h000;
			13355: dout = 12'h000;
			13356: dout = 12'h000;
			13357: dout = 12'h000;
			13358: dout = 12'h000;
			13359: dout = 12'h000;
			13360: dout = 12'h000;
			13361: dout = 12'h000;
			13362: dout = 12'h000;
			13363: dout = 12'h000;
			13364: dout = 12'h000;
			13365: dout = 12'h000;
			13366: dout = 12'h000;
			13367: dout = 12'h000;
			13368: dout = 12'h000;
			13369: dout = 12'h000;
			13370: dout = 12'h000;
			13371: dout = 12'h000;
			13372: dout = 12'haaa;
			13373: dout = 12'hfff;
			13374: dout = 12'h566;
			13375: dout = 12'h000;
			13376: dout = 12'h666;
			13377: dout = 12'hfff;
			13378: dout = 12'h000;
			13379: dout = 12'h000;
			13380: dout = 12'h000;
			13381: dout = 12'h000;
			13382: dout = 12'h000;
			13383: dout = 12'h000;
			13384: dout = 12'h000;
			13385: dout = 12'h000;
			13386: dout = 12'h000;
			13387: dout = 12'h000;
			13388: dout = 12'h000;
			13389: dout = 12'h000;
			13390: dout = 12'h000;
			13391: dout = 12'h000;
			13392: dout = 12'h000;
			13393: dout = 12'h000;
			13394: dout = 12'h000;
			13395: dout = 12'h000;
			13396: dout = 12'h000;
			13397: dout = 12'h000;
			13398: dout = 12'h000;
			13399: dout = 12'h555;
			13400: dout = 12'hfff;
			13401: dout = 12'habb;
			13402: dout = 12'hddd;
			13403: dout = 12'hfff;
			13404: dout = 12'hfff;
			13405: dout = 12'hfff;
			13406: dout = 12'haaa;
			13407: dout = 12'h000;
			13408: dout = 12'h000;
			13409: dout = 12'h000;
			13410: dout = 12'h000;
			13411: dout = 12'h000;
			13412: dout = 12'h000;
			13413: dout = 12'h333;
			13414: dout = 12'hfff;
			13415: dout = 12'hcdd;
			13416: dout = 12'habb;
			13417: dout = 12'habb;
			13418: dout = 12'hbbb;
			13419: dout = 12'h9aa;
			13420: dout = 12'hccc;
			13421: dout = 12'hfff;
			13422: dout = 12'hfff;
			13423: dout = 12'hfff;
			13424: dout = 12'h666;
			13425: dout = 12'h000;
			13426: dout = 12'h000;
			13427: dout = 12'h000;
			13428: dout = 12'h000;
			13429: dout = 12'h000;
			13430: dout = 12'h000;
			13431: dout = 12'h000;
			13432: dout = 12'h000;
			13433: dout = 12'h222;
			13434: dout = 12'hfff;
			13435: dout = 12'hfff;
			13436: dout = 12'hfff;
			13437: dout = 12'hfff;
			13438: dout = 12'hfff;
			13439: dout = 12'hfff;
			13440: dout = 12'hfff;
			13441: dout = 12'hfff;
			13442: dout = 12'hfff;
			13443: dout = 12'hfff;
			13444: dout = 12'hfff;
			13445: dout = 12'hfff;
			13446: dout = 12'h444;
			13447: dout = 12'h000;
			13448: dout = 12'h000;
			13449: dout = 12'h000;
			13450: dout = 12'h000;
			13451: dout = 12'h000;
			13452: dout = 12'h000;
			13453: dout = 12'h000;
			13454: dout = 12'h000;
			13455: dout = 12'h000;
			13456: dout = 12'h000;
			13457: dout = 12'h000;
			13458: dout = 12'h000;
			13459: dout = 12'h000;
			13460: dout = 12'h000;
			13461: dout = 12'h000;
			13462: dout = 12'h000;
			13463: dout = 12'h000;
			13464: dout = 12'h000;
			13465: dout = 12'h000;
			13466: dout = 12'h000;
			13467: dout = 12'h000;
			13468: dout = 12'h000;
			13469: dout = 12'h000;
			13470: dout = 12'h000;
			13471: dout = 12'h000;
			13472: dout = 12'h000;
			13473: dout = 12'h000;
			13474: dout = 12'h000;
			13475: dout = 12'h000;
			13476: dout = 12'h000;
			13477: dout = 12'h000;
			13478: dout = 12'h000;
			13479: dout = 12'h000;
			13480: dout = 12'h000;
			13481: dout = 12'h000;
			13482: dout = 12'h000;
			13483: dout = 12'h000;
			13484: dout = 12'h000;
			13485: dout = 12'h000;
			13486: dout = 12'h000;
			13487: dout = 12'h000;

			13488: dout = 12'h555;
			13489: dout = 12'hfff;
			13490: dout = 12'h100;
			13491: dout = 12'h600;
			13492: dout = 12'h500;
			13493: dout = 12'h400;
			13494: dout = 12'h400;
			13495: dout = 12'h300;
			13496: dout = 12'h000;
			13497: dout = 12'h000;
			13498: dout = 12'h000;
			13499: dout = 12'hfff;
			13500: dout = 12'hccc;
			13501: dout = 12'h000;
			13502: dout = 12'h000;
			13503: dout = 12'h000;
			13504: dout = 12'h000;
			13505: dout = 12'h000;
			13506: dout = 12'h000;
			13507: dout = 12'h000;
			13508: dout = 12'h000;
			13509: dout = 12'h000;
			13510: dout = 12'h000;
			13511: dout = 12'h000;
			13512: dout = 12'h000;
			13513: dout = 12'h000;
			13514: dout = 12'h000;
			13515: dout = 12'h000;
			13516: dout = 12'h000;
			13517: dout = 12'h000;
			13518: dout = 12'hfff;
			13519: dout = 12'h555;
			13520: dout = 12'hb10;
			13521: dout = 12'ha10;
			13522: dout = 12'h000;
			13523: dout = 12'hfff;
			13524: dout = 12'h444;
			13525: dout = 12'h000;
			13526: dout = 12'h000;
			13527: dout = 12'h000;
			13528: dout = 12'h000;
			13529: dout = 12'h000;
			13530: dout = 12'h000;
			13531: dout = 12'h000;
			13532: dout = 12'h000;
			13533: dout = 12'h000;
			13534: dout = 12'h000;
			13535: dout = 12'h000;
			13536: dout = 12'h000;
			13537: dout = 12'h000;
			13538: dout = 12'h000;
			13539: dout = 12'h000;
			13540: dout = 12'h000;
			13541: dout = 12'h000;
			13542: dout = 12'h000;
			13543: dout = 12'h000;
			13544: dout = 12'h111;
			13545: dout = 12'hfff;
			13546: dout = 12'h899;
			13547: dout = 12'h400;
			13548: dout = 12'h100;
			13549: dout = 12'h000;
			13550: dout = 12'h000;
			13551: dout = 12'h333;
			13552: dout = 12'hfff;
			13553: dout = 12'hccc;
			13554: dout = 12'h000;
			13555: dout = 12'h000;
			13556: dout = 12'h000;
			13557: dout = 12'h000;
			13558: dout = 12'h000;
			13559: dout = 12'hddd;
			13560: dout = 12'hbcc;
			13561: dout = 12'h300;
			13562: dout = 12'h600;
			13563: dout = 12'h400;
			13564: dout = 12'h400;
			13565: dout = 12'h300;
			13566: dout = 12'h100;
			13567: dout = 12'h000;
			13568: dout = 12'h000;
			13569: dout = 12'h777;
			13570: dout = 12'hfff;
			13571: dout = 12'h777;
			13572: dout = 12'h000;
			13573: dout = 12'h000;
			13574: dout = 12'h000;
			13575: dout = 12'h000;
			13576: dout = 12'h000;
			13577: dout = 12'h000;
			13578: dout = 12'h000;
			13579: dout = 12'hccc;
			13580: dout = 12'hccc;
			13581: dout = 12'h000;
			13582: dout = 12'h000;
			13583: dout = 12'h000;
			13584: dout = 12'h000;
			13585: dout = 12'haaa;
			13586: dout = 12'hddd;
			13587: dout = 12'h000;
			13588: dout = 12'h000;
			13589: dout = 12'h000;
			13590: dout = 12'h000;
			13591: dout = 12'haaa;
			13592: dout = 12'hfff;
			13593: dout = 12'h000;
			13594: dout = 12'h000;
			13595: dout = 12'h000;
			13596: dout = 12'h000;
			13597: dout = 12'h000;
			13598: dout = 12'h000;
			13599: dout = 12'h000;
			13600: dout = 12'h000;
			13601: dout = 12'h000;
			13602: dout = 12'h000;
			13603: dout = 12'h000;
			13604: dout = 12'h000;
			13605: dout = 12'h000;
			13606: dout = 12'h000;
			13607: dout = 12'h000;
			13608: dout = 12'h000;
			13609: dout = 12'h000;
			13610: dout = 12'h000;
			13611: dout = 12'h000;
			13612: dout = 12'h000;
			13613: dout = 12'h000;
			13614: dout = 12'h000;
			13615: dout = 12'h000;
			13616: dout = 12'h000;
			13617: dout = 12'h000;
			13618: dout = 12'h000;
			13619: dout = 12'h000;
			13620: dout = 12'h000;
			13621: dout = 12'h000;
			13622: dout = 12'h000;
			13623: dout = 12'h000;
			13624: dout = 12'h000;
			13625: dout = 12'h000;
			13626: dout = 12'h000;
			13627: dout = 12'h000;
			13628: dout = 12'h000;
			13629: dout = 12'h000;
			13630: dout = 12'h000;
			13631: dout = 12'h000;
			13632: dout = 12'h000;
			13633: dout = 12'h000;

			13634: dout = 12'h444;
			13635: dout = 12'hfff;
			13636: dout = 12'h200;
			13637: dout = 12'hc30;
			13638: dout = 12'he30;
			13639: dout = 12'hf40;
			13640: dout = 12'hc30;
			13641: dout = 12'hf40;
			13642: dout = 12'hf40;
			13643: dout = 12'hc30;
			13644: dout = 12'h000;
			13645: dout = 12'h455;
			13646: dout = 12'hfff;
			13647: dout = 12'hccc;
			13648: dout = 12'h000;
			13649: dout = 12'h000;
			13650: dout = 12'h000;
			13651: dout = 12'h000;
			13652: dout = 12'h000;
			13653: dout = 12'h000;
			13654: dout = 12'h000;
			13655: dout = 12'h000;
			13656: dout = 12'h000;
			13657: dout = 12'h000;
			13658: dout = 12'h000;
			13659: dout = 12'h000;
			13660: dout = 12'h000;
			13661: dout = 12'h000;
			13662: dout = 12'h000;
			13663: dout = 12'h000;
			13664: dout = 12'hfff;
			13665: dout = 12'h222;
			13666: dout = 12'hc20;
			13667: dout = 12'h710;
			13668: dout = 12'h000;
			13669: dout = 12'hfff;
			13670: dout = 12'hbbb;
			13671: dout = 12'h555;
			13672: dout = 12'h444;
			13673: dout = 12'h333;
			13674: dout = 12'h000;
			13675: dout = 12'h000;
			13676: dout = 12'h000;
			13677: dout = 12'h000;
			13678: dout = 12'h000;
			13679: dout = 12'h000;
			13680: dout = 12'h000;
			13681: dout = 12'h000;
			13682: dout = 12'h000;
			13683: dout = 12'h000;
			13684: dout = 12'h000;
			13685: dout = 12'h000;
			13686: dout = 12'h000;
			13687: dout = 12'h000;
			13688: dout = 12'h000;
			13689: dout = 12'h000;
			13690: dout = 12'hfff;
			13691: dout = 12'hddd;
			13692: dout = 12'h244;
			13693: dout = 12'hb20;
			13694: dout = 12'hd30;
			13695: dout = 12'hc30;
			13696: dout = 12'hd30;
			13697: dout = 12'h000;
			13698: dout = 12'h777;
			13699: dout = 12'hfff;
			13700: dout = 12'heee;
			13701: dout = 12'h000;
			13702: dout = 12'h000;
			13703: dout = 12'h000;
			13704: dout = 12'h000;
			13705: dout = 12'hccc;
			13706: dout = 12'habb;
			13707: dout = 12'h710;
			13708: dout = 12'hd30;
			13709: dout = 12'hf40;
			13710: dout = 12'hd30;
			13711: dout = 12'he30;
			13712: dout = 12'hf40;
			13713: dout = 12'hf40;
			13714: dout = 12'h610;
			13715: dout = 12'h000;
			13716: dout = 12'h788;
			13717: dout = 12'hfff;
			13718: dout = 12'h555;
			13719: dout = 12'h000;
			13720: dout = 12'h000;
			13721: dout = 12'h000;
			13722: dout = 12'h000;
			13723: dout = 12'h000;
			13724: dout = 12'h000;
			13725: dout = 12'hddd;
			13726: dout = 12'h899;
			13727: dout = 12'ha10;
			13728: dout = 12'he30;
			13729: dout = 12'hf30;
			13730: dout = 12'h710;
			13731: dout = 12'h001;
			13732: dout = 12'habb;
			13733: dout = 12'ha10;
			13734: dout = 12'he30;
			13735: dout = 12'hf30;
			13736: dout = 12'h710;
			13737: dout = 12'h000;
			13738: dout = 12'hfff;
			13739: dout = 12'h111;
			13740: dout = 12'h000;
			13741: dout = 12'h000;
			13742: dout = 12'h000;
			13743: dout = 12'h000;
			13744: dout = 12'h000;
			13745: dout = 12'h000;
			13746: dout = 12'h000;
			13747: dout = 12'h000;
			13748: dout = 12'h000;
			13749: dout = 12'h000;
			13750: dout = 12'h000;
			13751: dout = 12'h000;
			13752: dout = 12'h000;
			13753: dout = 12'h000;
			13754: dout = 12'h000;
			13755: dout = 12'h000;
			13756: dout = 12'h000;
			13757: dout = 12'h000;
			13758: dout = 12'h000;
			13759: dout = 12'h000;
			13760: dout = 12'h000;
			13761: dout = 12'h000;
			13762: dout = 12'h000;
			13763: dout = 12'h000;
			13764: dout = 12'h000;
			13765: dout = 12'h000;
			13766: dout = 12'h000;
			13767: dout = 12'h000;
			13768: dout = 12'h000;
			13769: dout = 12'h000;
			13770: dout = 12'h000;
			13771: dout = 12'h000;
			13772: dout = 12'h000;
			13773: dout = 12'h000;
			13774: dout = 12'h000;
			13775: dout = 12'h000;
			13776: dout = 12'h000;
			13777: dout = 12'h000;
			13778: dout = 12'h000;
			13779: dout = 12'h000;

			13780: dout = 12'h666;
			13781: dout = 12'hfff;
			13782: dout = 12'h300;
			13783: dout = 12'hd40;
			13784: dout = 12'h310;
			13785: dout = 12'h000;
			13786: dout = 12'h000;
			13787: dout = 12'h000;
			13788: dout = 12'h000;
			13789: dout = 12'h200;
			13790: dout = 12'hc30;
			13791: dout = 12'h400;
			13792: dout = 12'h333;
			13793: dout = 12'hfff;
			13794: dout = 12'heee;
			13795: dout = 12'heee;
			13796: dout = 12'hbbb;
			13797: dout = 12'hbbb;
			13798: dout = 12'hbbb;
			13799: dout = 12'hddd;
			13800: dout = 12'h666;
			13801: dout = 12'h999;
			13802: dout = 12'hfff;
			13803: dout = 12'hfff;
			13804: dout = 12'heee;
			13805: dout = 12'hfff;
			13806: dout = 12'hfff;
			13807: dout = 12'hccc;
			13808: dout = 12'hfff;
			13809: dout = 12'hfff;
			13810: dout = 12'hfff;
			13811: dout = 12'h777;
			13812: dout = 12'hc30;
			13813: dout = 12'h920;
			13814: dout = 12'h000;
			13815: dout = 12'hfff;
			13816: dout = 12'hfff;
			13817: dout = 12'hfff;
			13818: dout = 12'hfff;
			13819: dout = 12'hfff;
			13820: dout = 12'hfff;
			13821: dout = 12'h000;
			13822: dout = 12'h000;
			13823: dout = 12'h666;
			13824: dout = 12'h555;
			13825: dout = 12'h777;
			13826: dout = 12'h999;
			13827: dout = 12'haaa;
			13828: dout = 12'hfff;
			13829: dout = 12'hddd;
			13830: dout = 12'hccc;
			13831: dout = 12'haaa;
			13832: dout = 12'h000;
			13833: dout = 12'h000;
			13834: dout = 12'h000;
			13835: dout = 12'h999;
			13836: dout = 12'hfff;
			13837: dout = 12'h200;
			13838: dout = 12'h820;
			13839: dout = 12'ha30;
			13840: dout = 12'h920;
			13841: dout = 12'h920;
			13842: dout = 12'ha30;
			13843: dout = 12'hb30;
			13844: dout = 12'h200;
			13845: dout = 12'h233;
			13846: dout = 12'hfff;
			13847: dout = 12'h000;
			13848: dout = 12'h000;
			13849: dout = 12'h000;
			13850: dout = 12'h000;
			13851: dout = 12'hddd;
			13852: dout = 12'h9aa;
			13853: dout = 12'h810;
			13854: dout = 12'hc30;
			13855: dout = 12'h000;
			13856: dout = 12'h000;
			13857: dout = 12'h000;
			13858: dout = 12'h100;
			13859: dout = 12'h000;
			13860: dout = 12'h510;
			13861: dout = 12'hd30;
			13862: dout = 12'h000;
			13863: dout = 12'h999;
			13864: dout = 12'hfff;
			13865: dout = 12'hfff;
			13866: dout = 12'hfff;
			13867: dout = 12'hfff;
			13868: dout = 12'hfff;
			13869: dout = 12'hfff;
			13870: dout = 12'hfff;
			13871: dout = 12'hfff;
			13872: dout = 12'h899;
			13873: dout = 12'h400;
			13874: dout = 12'h820;
			13875: dout = 12'ha30;
			13876: dout = 12'h920;
			13877: dout = 12'h000;
			13878: dout = 12'habb;
			13879: dout = 12'h400;
			13880: dout = 12'h720;
			13881: dout = 12'ha30;
			13882: dout = 12'h920;
			13883: dout = 12'h000;
			13884: dout = 12'hfff;
			13885: dout = 12'h222;
			13886: dout = 12'haaa;
			13887: dout = 12'hfff;
			13888: dout = 12'hddd;
			13889: dout = 12'hbbb;
			13890: dout = 12'hbbb;
			13891: dout = 12'hccc;
			13892: dout = 12'hccc;
			13893: dout = 12'h444;
			13894: dout = 12'h000;
			13895: dout = 12'h333;
			13896: dout = 12'hddd;
			13897: dout = 12'hfff;
			13898: dout = 12'hbbb;
			13899: dout = 12'hbbb;
			13900: dout = 12'hbbb;
			13901: dout = 12'hddd;
			13902: dout = 12'h999;
			13903: dout = 12'h777;
			13904: dout = 12'hfff;
			13905: dout = 12'hfff;
			13906: dout = 12'hfff;
			13907: dout = 12'hfff;
			13908: dout = 12'hfff;
			13909: dout = 12'hfff;
			13910: dout = 12'hfff;
			13911: dout = 12'hfff;
			13912: dout = 12'hfff;
			13913: dout = 12'h111;
			13914: dout = 12'h000;
			13915: dout = 12'h444;
			13916: dout = 12'h555;
			13917: dout = 12'h555;
			13918: dout = 12'h999;
			13919: dout = 12'h999;
			13920: dout = 12'heee;
			13921: dout = 12'heee;
			13922: dout = 12'hccc;
			13923: dout = 12'hccc;
			13924: dout = 12'h333;
			13925: dout = 12'h000;

			13926: dout = 12'h888;
			13927: dout = 12'heef;
			13928: dout = 12'h200;
			13929: dout = 12'hf50;
			13930: dout = 12'h000;
			13931: dout = 12'h888;
			13932: dout = 12'hbbb;
			13933: dout = 12'hbbb;
			13934: dout = 12'hbbb;
			13935: dout = 12'h455;
			13936: dout = 12'hb30;
			13937: dout = 12'h720;
			13938: dout = 12'h000;
			13939: dout = 12'hfff;
			13940: dout = 12'h788;
			13941: dout = 12'h99a;
			13942: dout = 12'hbcc;
			13943: dout = 12'hccd;
			13944: dout = 12'hbbc;
			13945: dout = 12'haaa;
			13946: dout = 12'hfff;
			13947: dout = 12'hfff;
			13948: dout = 12'h566;
			13949: dout = 12'h889;
			13950: dout = 12'h899;
			13951: dout = 12'h889;
			13952: dout = 12'h999;
			13953: dout = 12'heff;
			13954: dout = 12'h556;
			13955: dout = 12'h334;
			13956: dout = 12'hfff;
			13957: dout = 12'h443;
			13958: dout = 12'hd40;
			13959: dout = 12'hb30;
			13960: dout = 12'h001;
			13961: dout = 12'h321;
			13962: dout = 12'h100;
			13963: dout = 12'h000;
			13964: dout = 12'h000;
			13965: dout = 12'h000;
			13966: dout = 12'heee;
			13967: dout = 12'hfff;
			13968: dout = 12'hfff;
			13969: dout = 12'hfff;
			13970: dout = 12'hfff;
			13971: dout = 12'hfff;
			13972: dout = 12'hdee;
			13973: dout = 12'hdee;
			13974: dout = 12'h788;
			13975: dout = 12'haab;
			13976: dout = 12'haaa;
			13977: dout = 12'hfff;
			13978: dout = 12'heee;
			13979: dout = 12'h000;
			13980: dout = 12'h000;
			13981: dout = 12'hddd;
			13982: dout = 12'h9aa;
			13983: dout = 12'h920;
			13984: dout = 12'hc40;
			13985: dout = 12'h000;
			13986: dout = 12'h000;
			13987: dout = 12'h000;
			13988: dout = 12'h000;
			13989: dout = 12'hf50;
			13990: dout = 12'h830;
			13991: dout = 12'h000;
			13992: dout = 12'hfff;
			13993: dout = 12'h333;
			13994: dout = 12'h000;
			13995: dout = 12'h000;
			13996: dout = 12'h000;
			13997: dout = 12'hfff;
			13998: dout = 12'h788;
			13999: dout = 12'h820;
			14000: dout = 12'hb40;
			14001: dout = 12'h000;
			14002: dout = 12'hccc;
			14003: dout = 12'hbbc;
			14004: dout = 12'habb;
			14005: dout = 12'hbbc;
			14006: dout = 12'h221;
			14007: dout = 12'he40;
			14008: dout = 12'h200;
			14009: dout = 12'h445;
			14010: dout = 12'heee;
			14011: dout = 12'h122;
			14012: dout = 12'h122;
			14013: dout = 12'h234;
			14014: dout = 12'h233;
			14015: dout = 12'h455;
			14016: dout = 12'h888;
			14017: dout = 12'hfff;
			14018: dout = 12'hfff;
			14019: dout = 12'h344;
			14020: dout = 12'h122;
			14021: dout = 12'hc40;
			14022: dout = 12'h820;
			14023: dout = 12'h000;
			14024: dout = 12'hfff;
			14025: dout = 12'h344;
			14026: dout = 12'h122;
			14027: dout = 12'hc40;
			14028: dout = 12'h820;
			14029: dout = 12'h000;
			14030: dout = 12'hfff;
			14031: dout = 12'hfff;
			14032: dout = 12'hfff;
			14033: dout = 12'h677;
			14034: dout = 12'habb;
			14035: dout = 12'hccc;
			14036: dout = 12'hccd;
			14037: dout = 12'habb;
			14038: dout = 12'hccc;
			14039: dout = 12'hfff;
			14040: dout = 12'h777;
			14041: dout = 12'hfff;
			14042: dout = 12'habb;
			14043: dout = 12'h788;
			14044: dout = 12'hbcc;
			14045: dout = 12'hccc;
			14046: dout = 12'hbcc;
			14047: dout = 12'h9aa;
			14048: dout = 12'hfff;
			14049: dout = 12'hfff;
			14050: dout = 12'h677;
			14051: dout = 12'h123;
			14052: dout = 12'h666;
			14053: dout = 12'hccc;
			14054: dout = 12'h122;
			14055: dout = 12'h233;
			14056: dout = 12'h344;
			14057: dout = 12'h223;
			14058: dout = 12'hccc;
			14059: dout = 12'hfff;
			14060: dout = 12'hbbb;
			14061: dout = 12'hfff;
			14062: dout = 12'hfff;
			14063: dout = 12'hfff;
			14064: dout = 12'heee;
			14065: dout = 12'heff;
			14066: dout = 12'h89a;
			14067: dout = 12'h899;
			14068: dout = 12'haab;
			14069: dout = 12'hccc;
			14070: dout = 12'hfff;
			14071: dout = 12'h111;

			14072: dout = 12'h999;
			14073: dout = 12'hfff;
			14074: dout = 12'h400;
			14075: dout = 12'hf60;
			14076: dout = 12'h000;
			14077: dout = 12'hccc;
			14078: dout = 12'hfff;
			14079: dout = 12'hfff;
			14080: dout = 12'hfff;
			14081: dout = 12'h99a;
			14082: dout = 12'hc40;
			14083: dout = 12'h310;
			14084: dout = 12'h233;
			14085: dout = 12'h99a;
			14086: dout = 12'h710;
			14087: dout = 12'h610;
			14088: dout = 12'h200;
			14089: dout = 12'h200;
			14090: dout = 12'h720;
			14091: dout = 12'h200;
			14092: dout = 12'h445;
			14093: dout = 12'h899;
			14094: dout = 12'h920;
			14095: dout = 12'h720;
			14096: dout = 12'h620;
			14097: dout = 12'h920;
			14098: dout = 12'h000;
			14099: dout = 12'h200;
			14100: dout = 12'ha30;
			14101: dout = 12'h000;
			14102: dout = 12'h888;
			14103: dout = 12'h333;
			14104: dout = 12'ha30;
			14105: dout = 12'h930;
			14106: dout = 12'h000;
			14107: dout = 12'h720;
			14108: dout = 12'hf60;
			14109: dout = 12'hf60;
			14110: dout = 12'he50;
			14111: dout = 12'h200;
			14112: dout = 12'h011;
			14113: dout = 12'hfff;
			14114: dout = 12'hfff;
			14115: dout = 12'h000;
			14116: dout = 12'h100;
			14117: dout = 12'h200;
			14118: dout = 12'h400;
			14119: dout = 12'h510;
			14120: dout = 12'h920;
			14121: dout = 12'h820;
			14122: dout = 12'h300;
			14123: dout = 12'h011;
			14124: dout = 12'hfff;
			14125: dout = 12'h111;
			14126: dout = 12'h000;
			14127: dout = 12'h999;
			14128: dout = 12'hdee;
			14129: dout = 12'h720;
			14130: dout = 12'ha40;
			14131: dout = 12'h000;
			14132: dout = 12'h433;
			14133: dout = 12'hf60;
			14134: dout = 12'hd50;
			14135: dout = 12'h000;
			14136: dout = 12'h000;
			14137: dout = 12'h555;
			14138: dout = 12'hfff;
			14139: dout = 12'h000;
			14140: dout = 12'h000;
			14141: dout = 12'h000;
			14142: dout = 12'h000;
			14143: dout = 12'hfff;
			14144: dout = 12'h899;
			14145: dout = 12'ha30;
			14146: dout = 12'h930;
			14147: dout = 12'h000;
			14148: dout = 12'hfff;
			14149: dout = 12'hfff;
			14150: dout = 12'hfff;
			14151: dout = 12'hfff;
			14152: dout = 12'h433;
			14153: dout = 12'he50;
			14154: dout = 12'h000;
			14155: dout = 12'h999;
			14156: dout = 12'h332;
			14157: dout = 12'he50;
			14158: dout = 12'he50;
			14159: dout = 12'ha30;
			14160: dout = 12'h930;
			14161: dout = 12'ha30;
			14162: dout = 12'h000;
			14163: dout = 12'hccc;
			14164: dout = 12'hfff;
			14165: dout = 12'hfff;
			14166: dout = 12'h433;
			14167: dout = 12'hd50;
			14168: dout = 12'h720;
			14169: dout = 12'h001;
			14170: dout = 12'hfff;
			14171: dout = 12'hfff;
			14172: dout = 12'h444;
			14173: dout = 12'hd50;
			14174: dout = 12'h730;
			14175: dout = 12'h000;
			14176: dout = 12'hfff;
			14177: dout = 12'hfff;
			14178: dout = 12'h222;
			14179: dout = 12'h930;
			14180: dout = 12'h510;
			14181: dout = 12'h000;
			14182: dout = 12'h400;
			14183: dout = 12'h820;
			14184: dout = 12'h000;
			14185: dout = 12'h999;
			14186: dout = 12'hfff;
			14187: dout = 12'heef;
			14188: dout = 12'h300;
			14189: dout = 12'h820;
			14190: dout = 12'h410;
			14191: dout = 12'h000;
			14192: dout = 12'h510;
			14193: dout = 12'h610;
			14194: dout = 12'h000;
			14195: dout = 12'hbbc;
			14196: dout = 12'h710;
			14197: dout = 12'he50;
			14198: dout = 12'h000;
			14199: dout = 12'h333;
			14200: dout = 12'hd40;
			14201: dout = 12'h720;
			14202: dout = 12'hd50;
			14203: dout = 12'h820;
			14204: dout = 12'h000;
			14205: dout = 12'hfff;
			14206: dout = 12'hfff;
			14207: dout = 12'h332;
			14208: dout = 12'h100;
			14209: dout = 12'h100;
			14210: dout = 12'h400;
			14211: dout = 12'h300;
			14212: dout = 12'h820;
			14213: dout = 12'h720;
			14214: dout = 12'h820;
			14215: dout = 12'h000;
			14216: dout = 12'hddd;
			14217: dout = 12'haaa;

			14218: dout = 12'h555;
			14219: dout = 12'hfff;
			14220: dout = 12'h400;
			14221: dout = 12'hf60;
			14222: dout = 12'h000;
			14223: dout = 12'h112;
			14224: dout = 12'h444;
			14225: dout = 12'h566;
			14226: dout = 12'h566;
			14227: dout = 12'h012;
			14228: dout = 12'hd50;
			14229: dout = 12'hc50;
			14230: dout = 12'h000;
			14231: dout = 12'h345;
			14232: dout = 12'hd50;
			14233: dout = 12'hf70;
			14234: dout = 12'hb50;
			14235: dout = 12'hd60;
			14236: dout = 12'hc50;
			14237: dout = 12'ha40;
			14238: dout = 12'h000;
			14239: dout = 12'h123;
			14240: dout = 12'hc50;
			14241: dout = 12'h410;
			14242: dout = 12'he60;
			14243: dout = 12'he60;
			14244: dout = 12'h000;
			14245: dout = 12'h630;
			14246: dout = 12'hd60;
			14247: dout = 12'ha40;
			14248: dout = 12'h000;
			14249: dout = 12'h222;
			14250: dout = 12'hc50;
			14251: dout = 12'hd50;
			14252: dout = 12'h100;
			14253: dout = 12'hc50;
			14254: dout = 12'ha40;
			14255: dout = 12'h830;
			14256: dout = 12'h620;
			14257: dout = 12'hc50;
			14258: dout = 12'h620;
			14259: dout = 12'h000;
			14260: dout = 12'h567;
			14261: dout = 12'hb40;
			14262: dout = 12'hf70;
			14263: dout = 12'hf70;
			14264: dout = 12'hf70;
			14265: dout = 12'hf70;
			14266: dout = 12'hf60;
			14267: dout = 12'hf70;
			14268: dout = 12'h830;
			14269: dout = 12'h011;
			14270: dout = 12'hfff;
			14271: dout = 12'h111;
			14272: dout = 12'h000;
			14273: dout = 12'h777;
			14274: dout = 12'hfff;
			14275: dout = 12'h200;
			14276: dout = 12'hf60;
			14277: dout = 12'h000;
			14278: dout = 12'h000;
			14279: dout = 12'hf70;
			14280: dout = 12'hb50;
			14281: dout = 12'h000;
			14282: dout = 12'h777;
			14283: dout = 12'hfff;
			14284: dout = 12'h888;
			14285: dout = 12'h000;
			14286: dout = 12'h000;
			14287: dout = 12'h000;
			14288: dout = 12'h000;
			14289: dout = 12'hddd;
			14290: dout = 12'h9ab;
			14291: dout = 12'h930;
			14292: dout = 12'hc50;
			14293: dout = 12'h000;
			14294: dout = 12'h334;
			14295: dout = 12'h444;
			14296: dout = 12'h667;
			14297: dout = 12'h556;
			14298: dout = 12'h110;
			14299: dout = 12'hf70;
			14300: dout = 12'h620;
			14301: dout = 12'h344;
			14302: dout = 12'h333;
			14303: dout = 12'hc50;
			14304: dout = 12'hd50;
			14305: dout = 12'he60;
			14306: dout = 12'hc50;
			14307: dout = 12'he60;
			14308: dout = 12'h730;
			14309: dout = 12'h000;
			14310: dout = 12'h000;
			14311: dout = 12'hfff;
			14312: dout = 12'h223;
			14313: dout = 12'he60;
			14314: dout = 12'h520;
			14315: dout = 12'h001;
			14316: dout = 12'hfff;
			14317: dout = 12'hfff;
			14318: dout = 12'h333;
			14319: dout = 12'he50;
			14320: dout = 12'h520;
			14321: dout = 12'h001;
			14322: dout = 12'hfff;
			14323: dout = 12'h89a;
			14324: dout = 12'h111;
			14325: dout = 12'hf70;
			14326: dout = 12'hf60;
			14327: dout = 12'ha40;
			14328: dout = 12'hd50;
			14329: dout = 12'hd60;
			14330: dout = 12'h520;
			14331: dout = 12'h001;
			14332: dout = 12'h777;
			14333: dout = 12'h678;
			14334: dout = 12'h620;
			14335: dout = 12'hf70;
			14336: dout = 12'hd60;
			14337: dout = 12'hc50;
			14338: dout = 12'hc50;
			14339: dout = 12'hf60;
			14340: dout = 12'h000;
			14341: dout = 12'h123;
			14342: dout = 12'h410;
			14343: dout = 12'hb50;
			14344: dout = 12'h000;
			14345: dout = 12'h000;
			14346: dout = 12'hc50;
			14347: dout = 12'hb50;
			14348: dout = 12'hb50;
			14349: dout = 12'hb50;
			14350: dout = 12'h000;
			14351: dout = 12'h233;
			14352: dout = 12'hbbc;
			14353: dout = 12'h300;
			14354: dout = 12'hf70;
			14355: dout = 12'hf70;
			14356: dout = 12'hf70;
			14357: dout = 12'hf70;
			14358: dout = 12'hf60;
			14359: dout = 12'hf70;
			14360: dout = 12'hf70;
			14361: dout = 12'h000;
			14362: dout = 12'hccc;
			14363: dout = 12'haaa;

			14364: dout = 12'h555;
			14365: dout = 12'hfff;
			14366: dout = 12'h410;
			14367: dout = 12'he70;
			14368: dout = 12'ha50;
			14369: dout = 12'hd60;
			14370: dout = 12'h520;
			14371: dout = 12'h200;
			14372: dout = 12'h310;
			14373: dout = 12'h730;
			14374: dout = 12'h000;
			14375: dout = 12'h000;
			14376: dout = 12'h630;
			14377: dout = 12'hb50;
			14378: dout = 12'h420;
			14379: dout = 12'h000;
			14380: dout = 12'h000;
			14381: dout = 12'h000;
			14382: dout = 12'h000;
			14383: dout = 12'h940;
			14384: dout = 12'he60;
			14385: dout = 12'h310;
			14386: dout = 12'h410;
			14387: dout = 12'h730;
			14388: dout = 12'h100;
			14389: dout = 12'h310;
			14390: dout = 12'hc60;
			14391: dout = 12'hc60;
			14392: dout = 12'h000;
			14393: dout = 12'ha50;
			14394: dout = 12'hf70;
			14395: dout = 12'h100;
			14396: dout = 12'hd60;
			14397: dout = 12'he70;
			14398: dout = 12'hf80;
			14399: dout = 12'h000;
			14400: dout = 12'h000;
			14401: dout = 12'h112;
			14402: dout = 12'h011;
			14403: dout = 12'h940;
			14404: dout = 12'hf70;
			14405: dout = 12'h310;
			14406: dout = 12'h940;
			14407: dout = 12'h000;
			14408: dout = 12'h000;
			14409: dout = 12'h000;
			14410: dout = 12'h100;
			14411: dout = 12'h100;
			14412: dout = 12'h310;
			14413: dout = 12'h100;
			14414: dout = 12'h000;
			14415: dout = 12'h444;
			14416: dout = 12'hfff;
			14417: dout = 12'h000;
			14418: dout = 12'h000;
			14419: dout = 12'h222;
			14420: dout = 12'hfff;
			14421: dout = 12'h455;
			14422: dout = 12'h000;
			14423: dout = 12'hf80;
			14424: dout = 12'hf70;
			14425: dout = 12'h000;
			14426: dout = 12'h000;
			14427: dout = 12'h333;
			14428: dout = 12'hfff;
			14429: dout = 12'hfff;
			14430: dout = 12'hfff;
			14431: dout = 12'heee;
			14432: dout = 12'h000;
			14433: dout = 12'h000;
			14434: dout = 12'h000;
			14435: dout = 12'hccc;
			14436: dout = 12'haab;
			14437: dout = 12'ha40;
			14438: dout = 12'hd60;
			14439: dout = 12'hb50;
			14440: dout = 12'hd60;
			14441: dout = 12'h310;
			14442: dout = 12'h200;
			14443: dout = 12'h410;
			14444: dout = 12'h630;
			14445: dout = 12'h000;
			14446: dout = 12'h000;
			14447: dout = 12'h666;
			14448: dout = 12'hfff;
			14449: dout = 12'h000;
			14450: dout = 12'h000;
			14451: dout = 12'h000;
			14452: dout = 12'h000;
			14453: dout = 12'h000;
			14454: dout = 12'he70;
			14455: dout = 12'hf70;
			14456: dout = 12'h000;
			14457: dout = 12'hddd;
			14458: dout = 12'h433;
			14459: dout = 12'hf70;
			14460: dout = 12'h520;
			14461: dout = 12'h223;
			14462: dout = 12'hfff;
			14463: dout = 12'hfff;
			14464: dout = 12'h321;
			14465: dout = 12'hf70;
			14466: dout = 12'h520;
			14467: dout = 12'h222;
			14468: dout = 12'h99a;
			14469: dout = 12'h720;
			14470: dout = 12'ha50;
			14471: dout = 12'h210;
			14472: dout = 12'h000;
			14473: dout = 12'h000;
			14474: dout = 12'h000;
			14475: dout = 12'h000;
			14476: dout = 12'hd60;
			14477: dout = 12'hc60;
			14478: dout = 12'h100;
			14479: dout = 12'ha40;
			14480: dout = 12'h830;
			14481: dout = 12'h100;
			14482: dout = 12'h000;
			14483: dout = 12'h000;
			14484: dout = 12'h000;
			14485: dout = 12'h310;
			14486: dout = 12'hf70;
			14487: dout = 12'h830;
			14488: dout = 12'h520;
			14489: dout = 12'hb50;
			14490: dout = 12'hf70;
			14491: dout = 12'hf70;
			14492: dout = 12'h000;
			14493: dout = 12'h000;
			14494: dout = 12'h000;
			14495: dout = 12'h730;
			14496: dout = 12'hf80;
			14497: dout = 12'h410;
			14498: dout = 12'h720;
			14499: dout = 12'h520;
			14500: dout = 12'h000;
			14501: dout = 12'h000;
			14502: dout = 12'h000;
			14503: dout = 12'h000;
			14504: dout = 12'h310;
			14505: dout = 12'h100;
			14506: dout = 12'h100;
			14507: dout = 12'h000;
			14508: dout = 12'hfff;
			14509: dout = 12'h666;

			14510: dout = 12'h666;
			14511: dout = 12'hfff;
			14512: dout = 12'h100;
			14513: dout = 12'he70;
			14514: dout = 12'h950;
			14515: dout = 12'h630;
			14516: dout = 12'he70;
			14517: dout = 12'h730;
			14518: dout = 12'hc60;
			14519: dout = 12'hc60;
			14520: dout = 12'h310;
			14521: dout = 12'h000;
			14522: dout = 12'h420;
			14523: dout = 12'hc60;
			14524: dout = 12'h000;
			14525: dout = 12'h888;
			14526: dout = 12'haaa;
			14527: dout = 12'hcdd;
			14528: dout = 12'hcdd;
			14529: dout = 12'h100;
			14530: dout = 12'hf80;
			14531: dout = 12'h520;
			14532: dout = 12'h740;
			14533: dout = 12'hf80;
			14534: dout = 12'h000;
			14535: dout = 12'h210;
			14536: dout = 12'hf70;
			14537: dout = 12'h940;
			14538: dout = 12'h000;
			14539: dout = 12'h730;
			14540: dout = 12'hf80;
			14541: dout = 12'h310;
			14542: dout = 12'he70;
			14543: dout = 12'h520;
			14544: dout = 12'h520;
			14545: dout = 12'h200;
			14546: dout = 12'h000;
			14547: dout = 12'hfff;
			14548: dout = 12'hfff;
			14549: dout = 12'h100;
			14550: dout = 12'h940;
			14551: dout = 12'h310;
			14552: dout = 12'hf90;
			14553: dout = 12'h630;
			14554: dout = 12'h001;
			14555: dout = 12'h445;
			14556: dout = 12'h000;
			14557: dout = 12'h000;
			14558: dout = 12'h000;
			14559: dout = 12'h889;
			14560: dout = 12'haaa;
			14561: dout = 12'hfff;
			14562: dout = 12'h888;
			14563: dout = 12'h000;
			14564: dout = 12'h000;
			14565: dout = 12'h555;
			14566: dout = 12'hfff;
			14567: dout = 12'h321;
			14568: dout = 12'h420;
			14569: dout = 12'h840;
			14570: dout = 12'hf80;
			14571: dout = 12'h630;
			14572: dout = 12'h000;
			14573: dout = 12'haaa;
			14574: dout = 12'h899;
			14575: dout = 12'h000;
			14576: dout = 12'h001;
			14577: dout = 12'hfff;
			14578: dout = 12'h888;
			14579: dout = 12'h000;
			14580: dout = 12'h000;
			14581: dout = 12'hddd;
			14582: dout = 12'h99a;
			14583: dout = 12'h620;
			14584: dout = 12'hd70;
			14585: dout = 12'h840;
			14586: dout = 12'h840;
			14587: dout = 12'hc60;
			14588: dout = 12'h840;
			14589: dout = 12'hc60;
			14590: dout = 12'ha50;
			14591: dout = 12'h210;
			14592: dout = 12'h011;
			14593: dout = 12'hfff;
			14594: dout = 12'h888;
			14595: dout = 12'h000;
			14596: dout = 12'h112;
			14597: dout = 12'h111;
			14598: dout = 12'h310;
			14599: dout = 12'h310;
			14600: dout = 12'h730;
			14601: dout = 12'he70;
			14602: dout = 12'h000;
			14603: dout = 12'h777;
			14604: dout = 12'h445;
			14605: dout = 12'hd60;
			14606: dout = 12'h310;
			14607: dout = 12'h455;
			14608: dout = 12'hfff;
			14609: dout = 12'hfff;
			14610: dout = 12'h344;
			14611: dout = 12'hd60;
			14612: dout = 12'h310;
			14613: dout = 12'h555;
			14614: dout = 12'h99a;
			14615: dout = 12'h830;
			14616: dout = 12'h840;
			14617: dout = 12'h000;
			14618: dout = 12'habb;
			14619: dout = 12'haaa;
			14620: dout = 12'hddd;
			14621: dout = 12'haab;
			14622: dout = 12'h410;
			14623: dout = 12'hf80;
			14624: dout = 12'h210;
			14625: dout = 12'hd60;
			14626: dout = 12'h200;
			14627: dout = 12'h344;
			14628: dout = 12'hbbb;
			14629: dout = 12'hbbb;
			14630: dout = 12'hddd;
			14631: dout = 12'h444;
			14632: dout = 12'hb50;
			14633: dout = 12'hc60;
			14634: dout = 12'h530;
			14635: dout = 12'hd70;
			14636: dout = 12'hd70;
			14637: dout = 12'hb60;
			14638: dout = 12'h000;
			14639: dout = 12'hfff;
			14640: dout = 12'hfff;
			14641: dout = 12'h410;
			14642: dout = 12'hf80;
			14643: dout = 12'h630;
			14644: dout = 12'he70;
			14645: dout = 12'he70;
			14646: dout = 12'h000;
			14647: dout = 12'h445;
			14648: dout = 12'h001;
			14649: dout = 12'h000;
			14650: dout = 12'h000;
			14651: dout = 12'h344;
			14652: dout = 12'hbbb;
			14653: dout = 12'heee;
			14654: dout = 12'hfff;
			14655: dout = 12'h000;

			14656: dout = 12'h888;
			14657: dout = 12'heff;
			14658: dout = 12'h310;
			14659: dout = 12'hf90;
			14660: dout = 12'h000;
			14661: dout = 12'h112;
			14662: dout = 12'h000;
			14663: dout = 12'h011;
			14664: dout = 12'h000;
			14665: dout = 12'h000;
			14666: dout = 12'he80;
			14667: dout = 12'h740;
			14668: dout = 12'h210;
			14669: dout = 12'hf90;
			14670: dout = 12'h000;
			14671: dout = 12'hccc;
			14672: dout = 12'hfff;
			14673: dout = 12'haaa;
			14674: dout = 12'hfff;
			14675: dout = 12'h321;
			14676: dout = 12'hf90;
			14677: dout = 12'h530;
			14678: dout = 12'h950;
			14679: dout = 12'hb60;
			14680: dout = 12'h000;
			14681: dout = 12'h000;
			14682: dout = 12'he80;
			14683: dout = 12'h740;
			14684: dout = 12'h000;
			14685: dout = 12'h420;
			14686: dout = 12'hf80;
			14687: dout = 12'h110;
			14688: dout = 12'hf80;
			14689: dout = 12'h320;
			14690: dout = 12'h112;
			14691: dout = 12'h888;
			14692: dout = 12'hddd;
			14693: dout = 12'hfff;
			14694: dout = 12'heff;
			14695: dout = 12'h630;
			14696: dout = 12'he80;
			14697: dout = 12'h000;
			14698: dout = 12'h000;
			14699: dout = 12'he80;
			14700: dout = 12'ha60;
			14701: dout = 12'h950;
			14702: dout = 12'hd70;
			14703: dout = 12'hc60;
			14704: dout = 12'h840;
			14705: dout = 12'h000;
			14706: dout = 12'hfff;
			14707: dout = 12'hfff;
			14708: dout = 12'h555;
			14709: dout = 12'h000;
			14710: dout = 12'h000;
			14711: dout = 12'haaa;
			14712: dout = 12'hccd;
			14713: dout = 12'h630;
			14714: dout = 12'hf90;
			14715: dout = 12'h000;
			14716: dout = 12'h000;
			14717: dout = 12'hf90;
			14718: dout = 12'hb60;
			14719: dout = 12'h000;
			14720: dout = 12'h520;
			14721: dout = 12'hfa0;
			14722: dout = 12'h000;
			14723: dout = 12'h899;
			14724: dout = 12'hfff;
			14725: dout = 12'h000;
			14726: dout = 12'h000;
			14727: dout = 12'hfff;
			14728: dout = 12'h788;
			14729: dout = 12'ha50;
			14730: dout = 12'hb60;
			14731: dout = 12'h000;
			14732: dout = 12'h112;
			14733: dout = 12'h000;
			14734: dout = 12'h112;
			14735: dout = 12'h000;
			14736: dout = 12'h210;
			14737: dout = 12'hf90;
			14738: dout = 12'h100;
			14739: dout = 12'h889;
			14740: dout = 12'h320;
			14741: dout = 12'hf80;
			14742: dout = 12'hf80;
			14743: dout = 12'hf80;
			14744: dout = 12'hf90;
			14745: dout = 12'hf90;
			14746: dout = 12'hf80;
			14747: dout = 12'hd70;
			14748: dout = 12'h000;
			14749: dout = 12'hddd;
			14750: dout = 12'h444;
			14751: dout = 12'hf80;
			14752: dout = 12'h630;
			14753: dout = 12'h112;
			14754: dout = 12'hfff;
			14755: dout = 12'hfff;
			14756: dout = 12'h444;
			14757: dout = 12'hf80;
			14758: dout = 12'h630;
			14759: dout = 12'h112;
			14760: dout = 12'hcdd;
			14761: dout = 12'h520;
			14762: dout = 12'hd70;
			14763: dout = 12'h000;
			14764: dout = 12'hfff;
			14765: dout = 12'heee;
			14766: dout = 12'hddd;
			14767: dout = 12'heef;
			14768: dout = 12'h520;
			14769: dout = 12'hf90;
			14770: dout = 12'h100;
			14771: dout = 12'hd70;
			14772: dout = 12'h520;
			14773: dout = 12'h334;
			14774: dout = 12'hfff;
			14775: dout = 12'haaa;
			14776: dout = 12'hfff;
			14777: dout = 12'h567;
			14778: dout = 12'hd70;
			14779: dout = 12'hc60;
			14780: dout = 12'h630;
			14781: dout = 12'h840;
			14782: dout = 12'h000;
			14783: dout = 12'h000;
			14784: dout = 12'h222;
			14785: dout = 12'hfff;
			14786: dout = 12'hfff;
			14787: dout = 12'h210;
			14788: dout = 12'ha50;
			14789: dout = 12'h740;
			14790: dout = 12'h000;
			14791: dout = 12'h950;
			14792: dout = 12'hd70;
			14793: dout = 12'h840;
			14794: dout = 12'hc60;
			14795: dout = 12'hb60;
			14796: dout = 12'hc70;
			14797: dout = 12'h000;
			14798: dout = 12'haaa;
			14799: dout = 12'hfff;
			14800: dout = 12'hccc;
			14801: dout = 12'h000;

			14802: dout = 12'h999;
			14803: dout = 12'hcdd;
			14804: dout = 12'h520;
			14805: dout = 12'hf90;
			14806: dout = 12'h000;
			14807: dout = 12'hbbb;
			14808: dout = 12'hfff;
			14809: dout = 12'hfff;
			14810: dout = 12'hfff;
			14811: dout = 12'h9ab;
			14812: dout = 12'ha60;
			14813: dout = 12'h630;
			14814: dout = 12'h530;
			14815: dout = 12'hc70;
			14816: dout = 12'h000;
			14817: dout = 12'haaa;
			14818: dout = 12'heee;
			14819: dout = 12'h444;
			14820: dout = 12'hfff;
			14821: dout = 12'h431;
			14822: dout = 12'hf90;
			14823: dout = 12'h530;
			14824: dout = 12'h850;
			14825: dout = 12'he80;
			14826: dout = 12'h000;
			14827: dout = 12'h110;
			14828: dout = 12'hf90;
			14829: dout = 12'h740;
			14830: dout = 12'h001;
			14831: dout = 12'h850;
			14832: dout = 12'hb60;
			14833: dout = 12'h210;
			14834: dout = 12'hf90;
			14835: dout = 12'h210;
			14836: dout = 12'h223;
			14837: dout = 12'hfff;
			14838: dout = 12'hfff;
			14839: dout = 12'hfff;
			14840: dout = 12'hdde;
			14841: dout = 12'h620;
			14842: dout = 12'hd70;
			14843: dout = 12'h000;
			14844: dout = 12'h678;
			14845: dout = 12'hb60;
			14846: dout = 12'hd80;
			14847: dout = 12'he80;
			14848: dout = 12'hf90;
			14849: dout = 12'he80;
			14850: dout = 12'he80;
			14851: dout = 12'h000;
			14852: dout = 12'h000;
			14853: dout = 12'h777;
			14854: dout = 12'hfff;
			14855: dout = 12'h000;
			14856: dout = 12'h000;
			14857: dout = 12'h888;
			14858: dout = 12'hfff;
			14859: dout = 12'h740;
			14860: dout = 12'hf90;
			14861: dout = 12'h000;
			14862: dout = 12'h012;
			14863: dout = 12'h740;
			14864: dout = 12'hd80;
			14865: dout = 12'h740;
			14866: dout = 12'h950;
			14867: dout = 12'hf90;
			14868: dout = 12'h630;
			14869: dout = 12'h222;
			14870: dout = 12'hfff;
			14871: dout = 12'h000;
			14872: dout = 12'h000;
			14873: dout = 12'hfff;
			14874: dout = 12'h567;
			14875: dout = 12'hb60;
			14876: dout = 12'hb60;
			14877: dout = 12'h000;
			14878: dout = 12'hfff;
			14879: dout = 12'hfff;
			14880: dout = 12'hfff;
			14881: dout = 12'hfff;
			14882: dout = 12'h334;
			14883: dout = 12'hf90;
			14884: dout = 12'h100;
			14885: dout = 12'h200;
			14886: dout = 12'h850;
			14887: dout = 12'ha60;
			14888: dout = 12'h520;
			14889: dout = 12'h320;
			14890: dout = 12'h210;
			14891: dout = 12'h000;
			14892: dout = 12'h320;
			14893: dout = 12'hf90;
			14894: dout = 12'h000;
			14895: dout = 12'hbcc;
			14896: dout = 12'h442;
			14897: dout = 12'hf90;
			14898: dout = 12'h520;
			14899: dout = 12'h001;
			14900: dout = 12'hfff;
			14901: dout = 12'hfff;
			14902: dout = 12'h432;
			14903: dout = 12'hf90;
			14904: dout = 12'h530;
			14905: dout = 12'h111;
			14906: dout = 12'habc;
			14907: dout = 12'h950;
			14908: dout = 12'ha60;
			14909: dout = 12'h000;
			14910: dout = 12'hfff;
			14911: dout = 12'haaa;
			14912: dout = 12'h999;
			14913: dout = 12'heff;
			14914: dout = 12'h530;
			14915: dout = 12'hf90;
			14916: dout = 12'h210;
			14917: dout = 12'he80;
			14918: dout = 12'h420;
			14919: dout = 12'h111;
			14920: dout = 12'hfff;
			14921: dout = 12'h444;
			14922: dout = 12'hfff;
			14923: dout = 12'h667;
			14924: dout = 12'hc70;
			14925: dout = 12'hc70;
			14926: dout = 12'h100;
			14927: dout = 12'hb60;
			14928: dout = 12'h000;
			14929: dout = 12'hfff;
			14930: dout = 12'hfff;
			14931: dout = 12'heee;
			14932: dout = 12'hfff;
			14933: dout = 12'h310;
			14934: dout = 12'hfa0;
			14935: dout = 12'h310;
			14936: dout = 12'h567;
			14937: dout = 12'h420;
			14938: dout = 12'hf90;
			14939: dout = 12'hf90;
			14940: dout = 12'hd80;
			14941: dout = 12'hfa0;
			14942: dout = 12'hf90;
			14943: dout = 12'h320;
			14944: dout = 12'h000;
			14945: dout = 12'h000;
			14946: dout = 12'hfff;
			14947: dout = 12'h666;

			14948: dout = 12'h777;
			14949: dout = 12'hfff;
			14950: dout = 12'h200;
			14951: dout = 12'hfa0;
			14952: dout = 12'h000;
			14953: dout = 12'haab;
			14954: dout = 12'hfff;
			14955: dout = 12'hfff;
			14956: dout = 12'hfff;
			14957: dout = 12'h445;
			14958: dout = 12'he90;
			14959: dout = 12'h640;
			14960: dout = 12'h640;
			14961: dout = 12'hfa0;
			14962: dout = 12'h000;
			14963: dout = 12'h667;
			14964: dout = 12'heef;
			14965: dout = 12'hfff;
			14966: dout = 12'hfff;
			14967: dout = 12'h321;
			14968: dout = 12'hfa0;
			14969: dout = 12'h420;
			14970: dout = 12'hb70;
			14971: dout = 12'h530;
			14972: dout = 12'h000;
			14973: dout = 12'h111;
			14974: dout = 12'he90;
			14975: dout = 12'h740;
			14976: dout = 12'h112;
			14977: dout = 12'h430;
			14978: dout = 12'h640;
			14979: dout = 12'h320;
			14980: dout = 12'hfb0;
			14981: dout = 12'h960;
			14982: dout = 12'h000;
			14983: dout = 12'h899;
			14984: dout = 12'heee;
			14985: dout = 12'h9aa;
			14986: dout = 12'h789;
			14987: dout = 12'h320;
			14988: dout = 12'he90;
			14989: dout = 12'h000;
			14990: dout = 12'hbcc;
			14991: dout = 12'h000;
			14992: dout = 12'h000;
			14993: dout = 12'h000;
			14994: dout = 12'h000;
			14995: dout = 12'h000;
			14996: dout = 12'h430;
			14997: dout = 12'hfb0;
			14998: dout = 12'ha60;
			14999: dout = 12'h001;
			15000: dout = 12'hfff;
			15001: dout = 12'h111;
			15002: dout = 12'h000;
			15003: dout = 12'haaa;
			15004: dout = 12'hcdd;
			15005: dout = 12'h420;
			15006: dout = 12'hfb0;
			15007: dout = 12'h000;
			15008: dout = 12'h788;
			15009: dout = 12'h123;
			15010: dout = 12'h210;
			15011: dout = 12'hfb0;
			15012: dout = 12'h530;
			15013: dout = 12'h000;
			15014: dout = 12'h000;
			15015: dout = 12'h999;
			15016: dout = 12'hfff;
			15017: dout = 12'h000;
			15018: dout = 12'h000;
			15019: dout = 12'hfff;
			15020: dout = 12'h889;
			15021: dout = 12'h850;
			15022: dout = 12'hb70;
			15023: dout = 12'h000;
			15024: dout = 12'hfff;
			15025: dout = 12'hfff;
			15026: dout = 12'hfff;
			15027: dout = 12'hfff;
			15028: dout = 12'h110;
			15029: dout = 12'hfb0;
			15030: dout = 12'h100;
			15031: dout = 12'hfa0;
			15032: dout = 12'hfa0;
			15033: dout = 12'h000;
			15034: dout = 12'h122;
			15035: dout = 12'h455;
			15036: dout = 12'h556;
			15037: dout = 12'h234;
			15038: dout = 12'hc70;
			15039: dout = 12'hfa0;
			15040: dout = 12'h000;
			15041: dout = 12'hccc;
			15042: dout = 12'h222;
			15043: dout = 12'hfa0;
			15044: dout = 12'h640;
			15045: dout = 12'h001;
			15046: dout = 12'hfff;
			15047: dout = 12'hfff;
			15048: dout = 12'h222;
			15049: dout = 12'hfa0;
			15050: dout = 12'h740;
			15051: dout = 12'h112;
			15052: dout = 12'h888;
			15053: dout = 12'h960;
			15054: dout = 12'hd80;
			15055: dout = 12'h000;
			15056: dout = 12'h99a;
			15057: dout = 12'hfff;
			15058: dout = 12'hfff;
			15059: dout = 12'heef;
			15060: dout = 12'h420;
			15061: dout = 12'hfa0;
			15062: dout = 12'h320;
			15063: dout = 12'he90;
			15064: dout = 12'h630;
			15065: dout = 12'h001;
			15066: dout = 12'hccd;
			15067: dout = 12'hfff;
			15068: dout = 12'hfff;
			15069: dout = 12'h667;
			15070: dout = 12'hc70;
			15071: dout = 12'hb70;
			15072: dout = 12'h640;
			15073: dout = 12'he90;
			15074: dout = 12'h000;
			15075: dout = 12'hfff;
			15076: dout = 12'h888;
			15077: dout = 12'h000;
			15078: dout = 12'hfff;
			15079: dout = 12'h210;
			15080: dout = 12'hd80;
			15081: dout = 12'h210;
			15082: dout = 12'h677;
			15083: dout = 12'h445;
			15084: dout = 12'h000;
			15085: dout = 12'h000;
			15086: dout = 12'h000;
			15087: dout = 12'h000;
			15088: dout = 12'h000;
			15089: dout = 12'hfa0;
			15090: dout = 12'hfc0;
			15091: dout = 12'h000;
			15092: dout = 12'hbbb;
			15093: dout = 12'haaa;

			15094: dout = 12'h555;
			15095: dout = 12'hfff;
			15096: dout = 12'h210;
			15097: dout = 12'hfb0;
			15098: dout = 12'h530;
			15099: dout = 12'h000;
			15100: dout = 12'h000;
			15101: dout = 12'h222;
			15102: dout = 12'h000;
			15103: dout = 12'h950;
			15104: dout = 12'h960;
			15105: dout = 12'h960;
			15106: dout = 12'h210;
			15107: dout = 12'ha70;
			15108: dout = 12'h850;
			15109: dout = 12'h530;
			15110: dout = 12'h100;
			15111: dout = 12'h000;
			15112: dout = 12'h000;
			15113: dout = 12'h430;
			15114: dout = 12'h960;
			15115: dout = 12'h210;
			15116: dout = 12'hd80;
			15117: dout = 12'h960;
			15118: dout = 12'h000;
			15119: dout = 12'h211;
			15120: dout = 12'hfa0;
			15121: dout = 12'h740;
			15122: dout = 12'h012;
			15123: dout = 12'h740;
			15124: dout = 12'hfb0;
			15125: dout = 12'h000;
			15126: dout = 12'h000;
			15127: dout = 12'h960;
			15128: dout = 12'hb70;
			15129: dout = 12'h000;
			15130: dout = 12'h100;
			15131: dout = 12'h210;
			15132: dout = 12'h850;
			15133: dout = 12'h850;
			15134: dout = 12'h000;
			15135: dout = 12'h000;
			15136: dout = 12'h100;
			15137: dout = 12'h012;
			15138: dout = 12'h112;
			15139: dout = 12'h011;
			15140: dout = 12'h000;
			15141: dout = 12'h000;
			15142: dout = 12'h850;
			15143: dout = 12'hd90;
			15144: dout = 12'h420;
			15145: dout = 12'h011;
			15146: dout = 12'hfff;
			15147: dout = 12'h000;
			15148: dout = 12'h000;
			15149: dout = 12'h333;
			15150: dout = 12'hfff;
			15151: dout = 12'h000;
			15152: dout = 12'h320;
			15153: dout = 12'hb70;
			15154: dout = 12'h420;
			15155: dout = 12'h100;
			15156: dout = 12'h530;
			15157: dout = 12'h750;
			15158: dout = 12'hea0;
			15159: dout = 12'hd90;
			15160: dout = 12'h210;
			15161: dout = 12'h666;
			15162: dout = 12'hfff;
			15163: dout = 12'h000;
			15164: dout = 12'h000;
			15165: dout = 12'hddd;
			15166: dout = 12'h9ab;
			15167: dout = 12'h950;
			15168: dout = 12'hfa0;
			15169: dout = 12'h320;
			15170: dout = 12'h000;
			15171: dout = 12'h001;
			15172: dout = 12'h111;
			15173: dout = 12'h000;
			15174: dout = 12'ha70;
			15175: dout = 12'ha70;
			15176: dout = 12'h530;
			15177: dout = 12'h320;
			15178: dout = 12'hc80;
			15179: dout = 12'ha70;
			15180: dout = 12'h000;
			15181: dout = 12'h320;
			15182: dout = 12'h420;
			15183: dout = 12'h530;
			15184: dout = 12'ha60;
			15185: dout = 12'he90;
			15186: dout = 12'h210;
			15187: dout = 12'h000;
			15188: dout = 12'h420;
			15189: dout = 12'ha60;
			15190: dout = 12'h960;
			15191: dout = 12'h000;
			15192: dout = 12'h000;
			15193: dout = 12'h000;
			15194: dout = 12'h420;
			15195: dout = 12'ha60;
			15196: dout = 12'h960;
			15197: dout = 12'h000;
			15198: dout = 12'h000;
			15199: dout = 12'h640;
			15200: dout = 12'hb70;
			15201: dout = 12'h640;
			15202: dout = 12'h420;
			15203: dout = 12'h000;
			15204: dout = 12'h000;
			15205: dout = 12'h000;
			15206: dout = 12'h640;
			15207: dout = 12'h960;
			15208: dout = 12'h000;
			15209: dout = 12'h960;
			15210: dout = 12'ha60;
			15211: dout = 12'h530;
			15212: dout = 12'h210;
			15213: dout = 12'h000;
			15214: dout = 12'h000;
			15215: dout = 12'h100;
			15216: dout = 12'h850;
			15217: dout = 12'h640;
			15218: dout = 12'h750;
			15219: dout = 12'hc80;
			15220: dout = 12'h000;
			15221: dout = 12'h999;
			15222: dout = 12'hddd;
			15223: dout = 12'h444;
			15224: dout = 12'hfff;
			15225: dout = 12'h420;
			15226: dout = 12'hfb0;
			15227: dout = 12'h000;
			15228: dout = 12'h320;
			15229: dout = 12'h000;
			15230: dout = 12'h334;
			15231: dout = 12'h001;
			15232: dout = 12'h000;
			15233: dout = 12'h000;
			15234: dout = 12'h110;
			15235: dout = 12'hd90;
			15236: dout = 12'hb70;
			15237: dout = 12'h000;
			15238: dout = 12'hfff;
			15239: dout = 12'h888;

			15240: dout = 12'h666;
			15241: dout = 12'hfff;
			15242: dout = 12'h310;
			15243: dout = 12'hfb0;
			15244: dout = 12'hfa0;
			15245: dout = 12'hea0;
			15246: dout = 12'hb80;
			15247: dout = 12'hfb0;
			15248: dout = 12'hfa0;
			15249: dout = 12'h960;
			15250: dout = 12'h000;
			15251: dout = 12'h001;
			15252: dout = 12'h333;
			15253: dout = 12'h001;
			15254: dout = 12'hfc0;
			15255: dout = 12'hc80;
			15256: dout = 12'hfb0;
			15257: dout = 12'hc80;
			15258: dout = 12'hfb0;
			15259: dout = 12'hc90;
			15260: dout = 12'h000;
			15261: dout = 12'h111;
			15262: dout = 12'hea0;
			15263: dout = 12'hfa0;
			15264: dout = 12'h000;
			15265: dout = 12'h000;
			15266: dout = 12'hfb0;
			15267: dout = 12'ha70;
			15268: dout = 12'h000;
			15269: dout = 12'hb80;
			15270: dout = 12'hb80;
			15271: dout = 12'h100;
			15272: dout = 12'h667;
			15273: dout = 12'h310;
			15274: dout = 12'hfc0;
			15275: dout = 12'hc80;
			15276: dout = 12'hfc0;
			15277: dout = 12'hfb0;
			15278: dout = 12'hfd0;
			15279: dout = 12'h320;
			15280: dout = 12'h112;
			15281: dout = 12'h640;
			15282: dout = 12'hfc0;
			15283: dout = 12'hfb0;
			15284: dout = 12'hea0;
			15285: dout = 12'hfb0;
			15286: dout = 12'hfa0;
			15287: dout = 12'hfb0;
			15288: dout = 12'hd90;
			15289: dout = 12'h000;
			15290: dout = 12'h000;
			15291: dout = 12'hddd;
			15292: dout = 12'hfff;
			15293: dout = 12'h000;
			15294: dout = 12'h000;
			15295: dout = 12'h000;
			15296: dout = 12'hfff;
			15297: dout = 12'hfff;
			15298: dout = 12'h112;
			15299: dout = 12'hfc0;
			15300: dout = 12'hfb0;
			15301: dout = 12'hfc0;
			15302: dout = 12'hea0;
			15303: dout = 12'h000;
			15304: dout = 12'h210;
			15305: dout = 12'hfd0;
			15306: dout = 12'h420;
			15307: dout = 12'h566;
			15308: dout = 12'hfff;
			15309: dout = 12'h000;
			15310: dout = 12'h000;
			15311: dout = 12'heee;
			15312: dout = 12'h899;
			15313: dout = 12'h960;
			15314: dout = 12'hea0;
			15315: dout = 12'hfb0;
			15316: dout = 12'hd90;
			15317: dout = 12'hd90;
			15318: dout = 12'hfa0;
			15319: dout = 12'hea0;
			15320: dout = 12'h530;
			15321: dout = 12'h000;
			15322: dout = 12'h000;
			15323: dout = 12'h556;
			15324: dout = 12'h430;
			15325: dout = 12'hb80;
			15326: dout = 12'hfc0;
			15327: dout = 12'hfc0;
			15328: dout = 12'hfc0;
			15329: dout = 12'hfc0;
			15330: dout = 12'hfb0;
			15331: dout = 12'hfc0;
			15332: dout = 12'h210;
			15333: dout = 12'hfa0;
			15334: dout = 12'hea0;
			15335: dout = 12'h640;
			15336: dout = 12'hfb0;
			15337: dout = 12'hfd0;
			15338: dout = 12'h960;
			15339: dout = 12'hea0;
			15340: dout = 12'hea0;
			15341: dout = 12'h640;
			15342: dout = 12'hfb0;
			15343: dout = 12'hfc0;
			15344: dout = 12'ha70;
			15345: dout = 12'h000;
			15346: dout = 12'h320;
			15347: dout = 12'hfc0;
			15348: dout = 12'hb80;
			15349: dout = 12'hfb0;
			15350: dout = 12'hd90;
			15351: dout = 12'hfc0;
			15352: dout = 12'h750;
			15353: dout = 12'h000;
			15354: dout = 12'h444;
			15355: dout = 12'h123;
			15356: dout = 12'ha70;
			15357: dout = 12'hfa0;
			15358: dout = 12'hea0;
			15359: dout = 12'hc90;
			15360: dout = 12'hfa0;
			15361: dout = 12'hfd0;
			15362: dout = 12'h000;
			15363: dout = 12'h001;
			15364: dout = 12'hb80;
			15365: dout = 12'hfd0;
			15366: dout = 12'h000;
			15367: dout = 12'h999;
			15368: dout = 12'hccc;
			15369: dout = 12'h999;
			15370: dout = 12'hccd;
			15371: dout = 12'h750;
			15372: dout = 12'hfc0;
			15373: dout = 12'h210;
			15374: dout = 12'hfb0;
			15375: dout = 12'hfc0;
			15376: dout = 12'hea0;
			15377: dout = 12'hfb0;
			15378: dout = 12'hfb0;
			15379: dout = 12'hfb0;
			15380: dout = 12'hfb0;
			15381: dout = 12'h220;
			15382: dout = 12'h000;
			15383: dout = 12'h666;
			15384: dout = 12'hfff;
			15385: dout = 12'h333;

			15386: dout = 12'h555;
			15387: dout = 12'hfff;
			15388: dout = 12'h000;
			15389: dout = 12'h210;
			15390: dout = 12'h430;
			15391: dout = 12'h640;
			15392: dout = 12'h530;
			15393: dout = 12'h000;
			15394: dout = 12'h320;
			15395: dout = 12'h640;
			15396: dout = 12'h000;
			15397: dout = 12'heee;
			15398: dout = 12'hfff;
			15399: dout = 12'h332;
			15400: dout = 12'hc80;
			15401: dout = 12'h860;
			15402: dout = 12'h750;
			15403: dout = 12'h750;
			15404: dout = 12'hb80;
			15405: dout = 12'h960;
			15406: dout = 12'h000;
			15407: dout = 12'h445;
			15408: dout = 12'h740;
			15409: dout = 12'ha70;
			15410: dout = 12'h000;
			15411: dout = 12'h111;
			15412: dout = 12'h860;
			15413: dout = 12'h430;
			15414: dout = 12'h000;
			15415: dout = 12'h640;
			15416: dout = 12'h860;
			15417: dout = 12'h000;
			15418: dout = 12'h888;
			15419: dout = 12'h556;
			15420: dout = 12'h210;
			15421: dout = 12'h000;
			15422: dout = 12'h000;
			15423: dout = 12'h000;
			15424: dout = 12'h000;
			15425: dout = 12'h000;
			15426: dout = 12'hccd;
			15427: dout = 12'h320;
			15428: dout = 12'ha70;
			15429: dout = 12'h960;
			15430: dout = 12'ha70;
			15431: dout = 12'ha70;
			15432: dout = 12'ha70;
			15433: dout = 12'ha70;
			15434: dout = 12'h750;
			15435: dout = 12'h000;
			15436: dout = 12'hfff;
			15437: dout = 12'hfff;
			15438: dout = 12'h111;
			15439: dout = 12'h000;
			15440: dout = 12'h000;
			15441: dout = 12'h000;
			15442: dout = 12'h000;
			15443: dout = 12'hfff;
			15444: dout = 12'h888;
			15445: dout = 12'h000;
			15446: dout = 12'h430;
			15447: dout = 12'h320;
			15448: dout = 12'h110;
			15449: dout = 12'h000;
			15450: dout = 12'h333;
			15451: dout = 12'h100;
			15452: dout = 12'h000;
			15453: dout = 12'h778;
			15454: dout = 12'hfff;
			15455: dout = 12'h000;
			15456: dout = 12'h000;
			15457: dout = 12'hddd;
			15458: dout = 12'haaa;
			15459: dout = 12'h310;
			15460: dout = 12'h210;
			15461: dout = 12'h430;
			15462: dout = 12'h640;
			15463: dout = 12'h420;
			15464: dout = 12'h100;
			15465: dout = 12'h320;
			15466: dout = 12'h430;
			15467: dout = 12'h000;
			15468: dout = 12'hfff;
			15469: dout = 12'hfff;
			15470: dout = 12'h222;
			15471: dout = 12'h430;
			15472: dout = 12'h320;
			15473: dout = 12'h000;
			15474: dout = 12'h110;
			15475: dout = 12'h000;
			15476: dout = 12'h000;
			15477: dout = 12'h320;
			15478: dout = 12'h000;
			15479: dout = 12'hc80;
			15480: dout = 12'hb80;
			15481: dout = 12'h640;
			15482: dout = 12'h640;
			15483: dout = 12'h530;
			15484: dout = 12'h320;
			15485: dout = 12'hb80;
			15486: dout = 12'hb80;
			15487: dout = 12'h640;
			15488: dout = 12'h640;
			15489: dout = 12'h540;
			15490: dout = 12'h320;
			15491: dout = 12'h000;
			15492: dout = 12'h541;
			15493: dout = 12'hb80;
			15494: dout = 12'h750;
			15495: dout = 12'h640;
			15496: dout = 12'h960;
			15497: dout = 12'hc80;
			15498: dout = 12'h430;
			15499: dout = 12'h112;
			15500: dout = 12'hfff;
			15501: dout = 12'hbbc;
			15502: dout = 12'h750;
			15503: dout = 12'ha70;
			15504: dout = 12'h750;
			15505: dout = 12'h640;
			15506: dout = 12'ha70;
			15507: dout = 12'hc90;
			15508: dout = 12'h000;
			15509: dout = 12'h455;
			15510: dout = 12'h530;
			15511: dout = 12'h860;
			15512: dout = 12'h000;
			15513: dout = 12'hbbb;
			15514: dout = 12'hccc;
			15515: dout = 12'haaa;
			15516: dout = 12'hbbb;
			15517: dout = 12'h320;
			15518: dout = 12'hb80;
			15519: dout = 12'h000;
			15520: dout = 12'h970;
			15521: dout = 12'h860;
			15522: dout = 12'ha70;
			15523: dout = 12'ha70;
			15524: dout = 12'ha70;
			15525: dout = 12'ha70;
			15526: dout = 12'ha70;
			15527: dout = 12'h000;
			15528: dout = 12'haaa;
			15529: dout = 12'hfff;
			15530: dout = 12'h777;
			15531: dout = 12'h000;

			15532: dout = 12'h111;
			15533: dout = 12'hfff;
			15534: dout = 12'h899;
			15535: dout = 12'h777;
			15536: dout = 12'h455;
			15537: dout = 12'h444;
			15538: dout = 12'h445;
			15539: dout = 12'haaa;
			15540: dout = 12'haaa;
			15541: dout = 12'h444;
			15542: dout = 12'h999;
			15543: dout = 12'hfff;
			15544: dout = 12'hfff;
			15545: dout = 12'hccc;
			15546: dout = 12'h001;
			15547: dout = 12'h223;
			15548: dout = 12'h334;
			15549: dout = 12'h445;
			15550: dout = 12'h123;
			15551: dout = 12'h001;
			15552: dout = 12'h666;
			15553: dout = 12'hfff;
			15554: dout = 12'h333;
			15555: dout = 12'h223;
			15556: dout = 12'h777;
			15557: dout = 12'hfff;
			15558: dout = 12'h223;
			15559: dout = 12'h444;
			15560: dout = 12'hccc;
			15561: dout = 12'h344;
			15562: dout = 12'h233;
			15563: dout = 12'h333;
			15564: dout = 12'heee;
			15565: dout = 12'hfff;
			15566: dout = 12'h666;
			15567: dout = 12'h999;
			15568: dout = 12'hfff;
			15569: dout = 12'hccc;
			15570: dout = 12'hfff;
			15571: dout = 12'heee;
			15572: dout = 12'hfff;
			15573: dout = 12'h888;
			15574: dout = 12'h122;
			15575: dout = 12'h223;
			15576: dout = 12'h223;
			15577: dout = 12'h223;
			15578: dout = 12'h223;
			15579: dout = 12'h223;
			15580: dout = 12'h223;
			15581: dout = 12'h999;
			15582: dout = 12'hfff;
			15583: dout = 12'h000;
			15584: dout = 12'h000;
			15585: dout = 12'h000;
			15586: dout = 12'h000;
			15587: dout = 12'h000;
			15588: dout = 12'h000;
			15589: dout = 12'h666;
			15590: dout = 12'hfff;
			15591: dout = 12'heee;
			15592: dout = 12'h445;
			15593: dout = 12'h667;
			15594: dout = 12'h556;
			15595: dout = 12'heee;
			15596: dout = 12'hfff;
			15597: dout = 12'hbbb;
			15598: dout = 12'hbbb;
			15599: dout = 12'hfff;
			15600: dout = 12'h666;
			15601: dout = 12'h000;
			15602: dout = 12'h000;
			15603: dout = 12'h888;
			15604: dout = 12'hfff;
			15605: dout = 12'h667;
			15606: dout = 12'h777;
			15607: dout = 12'h444;
			15608: dout = 12'h445;
			15609: dout = 12'h556;
			15610: dout = 12'hbbb;
			15611: dout = 12'h899;
			15612: dout = 12'h334;
			15613: dout = 12'hddd;
			15614: dout = 12'hfff;
			15615: dout = 12'hbbb;
			15616: dout = 12'hfff;
			15617: dout = 12'h444;
			15618: dout = 12'h999;
			15619: dout = 12'h999;
			15620: dout = 12'h666;
			15621: dout = 12'heee;
			15622: dout = 12'hbbb;
			15623: dout = 12'h444;
			15624: dout = 12'h999;
			15625: dout = 12'h011;
			15626: dout = 12'h001;
			15627: dout = 12'h333;
			15628: dout = 12'h334;
			15629: dout = 12'h445;
			15630: dout = 12'h444;
			15631: dout = 12'h112;
			15632: dout = 12'h001;
			15633: dout = 12'h333;
			15634: dout = 12'h334;
			15635: dout = 12'h445;
			15636: dout = 12'h333;
			15637: dout = 12'hbbb;
			15638: dout = 12'h788;
			15639: dout = 12'h012;
			15640: dout = 12'h223;
			15641: dout = 12'h445;
			15642: dout = 12'h334;
			15643: dout = 12'h123;
			15644: dout = 12'h001;
			15645: dout = 12'hbbb;
			15646: dout = 12'hfff;
			15647: dout = 12'hfff;
			15648: dout = 12'h122;
			15649: dout = 12'h112;
			15650: dout = 12'h334;
			15651: dout = 12'h455;
			15652: dout = 12'h223;
			15653: dout = 12'h012;
			15654: dout = 12'h222;
			15655: dout = 12'hfff;
			15656: dout = 12'h555;
			15657: dout = 12'h334;
			15658: dout = 12'h777;
			15659: dout = 12'hfff;
			15660: dout = 12'h444;
			15661: dout = 12'h777;
			15662: dout = 12'hfff;
			15663: dout = 12'h555;
			15664: dout = 12'h223;
			15665: dout = 12'h445;
			15666: dout = 12'h223;
			15667: dout = 12'h223;
			15668: dout = 12'h223;
			15669: dout = 12'h223;
			15670: dout = 12'h223;
			15671: dout = 12'h223;
			15672: dout = 12'h223;
			15673: dout = 12'h444;
			15674: dout = 12'hfff;
			15675: dout = 12'h999;
			15676: dout = 12'h000;
			15677: dout = 12'h000;

			15678: dout = 12'h000;
			15679: dout = 12'h555;
			15680: dout = 12'hfff;
			15681: dout = 12'hfff;
			15682: dout = 12'hfff;
			15683: dout = 12'hfff;
			15684: dout = 12'hfff;
			15685: dout = 12'heee;
			15686: dout = 12'hddd;
			15687: dout = 12'hfff;
			15688: dout = 12'hfff;
			15689: dout = 12'h544;
			15690: dout = 12'h111;
			15691: dout = 12'hfff;
			15692: dout = 12'hfff;
			15693: dout = 12'hfff;
			15694: dout = 12'hfff;
			15695: dout = 12'hfff;
			15696: dout = 12'hfff;
			15697: dout = 12'hfff;
			15698: dout = 12'hfff;
			15699: dout = 12'heee;
			15700: dout = 12'hfff;
			15701: dout = 12'hfff;
			15702: dout = 12'hfff;
			15703: dout = 12'heee;
			15704: dout = 12'hfff;
			15705: dout = 12'hfff;
			15706: dout = 12'heee;
			15707: dout = 12'hfff;
			15708: dout = 12'hfff;
			15709: dout = 12'hfff;
			15710: dout = 12'hddd;
			15711: dout = 12'h888;
			15712: dout = 12'hfff;
			15713: dout = 12'hfff;
			15714: dout = 12'h888;
			15715: dout = 12'hccc;
			15716: dout = 12'h999;
			15717: dout = 12'haaa;
			15718: dout = 12'h666;
			15719: dout = 12'hfff;
			15720: dout = 12'hfff;
			15721: dout = 12'hfff;
			15722: dout = 12'hfff;
			15723: dout = 12'hfff;
			15724: dout = 12'hfff;
			15725: dout = 12'hfff;
			15726: dout = 12'hfff;
			15727: dout = 12'hfff;
			15728: dout = 12'h555;
			15729: dout = 12'h000;
			15730: dout = 12'h000;
			15731: dout = 12'h000;
			15732: dout = 12'h000;
			15733: dout = 12'h000;
			15734: dout = 12'h000;
			15735: dout = 12'h000;
			15736: dout = 12'h333;
			15737: dout = 12'hccc;
			15738: dout = 12'hfff;
			15739: dout = 12'hfff;
			15740: dout = 12'hfff;
			15741: dout = 12'hbbb;
			15742: dout = 12'h666;
			15743: dout = 12'hccc;
			15744: dout = 12'hddd;
			15745: dout = 12'h555;
			15746: dout = 12'h000;
			15747: dout = 12'h000;
			15748: dout = 12'h000;
			15749: dout = 12'h000;
			15750: dout = 12'haaa;
			15751: dout = 12'hfff;
			15752: dout = 12'hfff;
			15753: dout = 12'hfff;
			15754: dout = 12'hfff;
			15755: dout = 12'hfff;
			15756: dout = 12'hccc;
			15757: dout = 12'hfff;
			15758: dout = 12'hfff;
			15759: dout = 12'hddd;
			15760: dout = 12'h111;
			15761: dout = 12'h000;
			15762: dout = 12'hbbb;
			15763: dout = 12'hfff;
			15764: dout = 12'hfff;
			15765: dout = 12'heee;
			15766: dout = 12'hfff;
			15767: dout = 12'hccc;
			15768: dout = 12'hddd;
			15769: dout = 12'hfff;
			15770: dout = 12'hfff;
			15771: dout = 12'hfff;
			15772: dout = 12'hfff;
			15773: dout = 12'hfff;
			15774: dout = 12'hfff;
			15775: dout = 12'hfff;
			15776: dout = 12'hfff;
			15777: dout = 12'hfff;
			15778: dout = 12'hfff;
			15779: dout = 12'hfff;
			15780: dout = 12'hfff;
			15781: dout = 12'hfff;
			15782: dout = 12'hfff;
			15783: dout = 12'hfff;
			15784: dout = 12'hfff;
			15785: dout = 12'hfff;
			15786: dout = 12'hfff;
			15787: dout = 12'hfff;
			15788: dout = 12'hfff;
			15789: dout = 12'hfff;
			15790: dout = 12'hfff;
			15791: dout = 12'hfff;
			15792: dout = 12'h333;
			15793: dout = 12'hccc;
			15794: dout = 12'hfff;
			15795: dout = 12'hfff;
			15796: dout = 12'hfff;
			15797: dout = 12'hfff;
			15798: dout = 12'hfff;
			15799: dout = 12'hfff;
			15800: dout = 12'hfff;
			15801: dout = 12'heee;
			15802: dout = 12'hfff;
			15803: dout = 12'hfff;
			15804: dout = 12'hfff;
			15805: dout = 12'h777;
			15806: dout = 12'h000;
			15807: dout = 12'h000;
			15808: dout = 12'h999;
			15809: dout = 12'hfff;
			15810: dout = 12'hfff;
			15811: dout = 12'hfff;
			15812: dout = 12'hfff;
			15813: dout = 12'hfff;
			15814: dout = 12'hfff;
			15815: dout = 12'hfff;
			15816: dout = 12'hfff;
			15817: dout = 12'hfff;
			15818: dout = 12'hfff;
			15819: dout = 12'hfff;
			15820: dout = 12'hbbb;
			15821: dout = 12'h000;
			15822: dout = 12'h000;
			15823: dout = 12'h000;

			15824: dout = 12'h000;
			15825: dout = 12'h000;
			15826: dout = 12'h000;
			15827: dout = 12'h000;
			15828: dout = 12'h000;
			15829: dout = 12'h000;
			15830: dout = 12'h000;
			15831: dout = 12'h000;
			15832: dout = 12'h000;
			15833: dout = 12'h000;
			15834: dout = 12'h000;
			15835: dout = 12'h000;
			15836: dout = 12'h000;
			15837: dout = 12'h000;
			15838: dout = 12'h000;
			15839: dout = 12'h000;
			15840: dout = 12'h000;
			15841: dout = 12'h000;
			15842: dout = 12'h000;
			15843: dout = 12'h000;
			15844: dout = 12'h000;
			15845: dout = 12'h000;
			15846: dout = 12'h000;
			15847: dout = 12'h000;
			15848: dout = 12'h000;
			15849: dout = 12'h000;
			15850: dout = 12'h000;
			15851: dout = 12'h000;
			15852: dout = 12'h000;
			15853: dout = 12'h000;
			15854: dout = 12'h000;
			15855: dout = 12'h000;
			15856: dout = 12'h000;
			15857: dout = 12'h000;
			15858: dout = 12'h000;
			15859: dout = 12'h000;
			15860: dout = 12'h000;
			15861: dout = 12'h000;
			15862: dout = 12'h000;
			15863: dout = 12'h000;
			15864: dout = 12'h000;
			15865: dout = 12'h000;
			15866: dout = 12'h000;
			15867: dout = 12'h000;
			15868: dout = 12'h000;
			15869: dout = 12'h000;
			15870: dout = 12'h000;
			15871: dout = 12'h000;
			15872: dout = 12'h000;
			15873: dout = 12'h000;
			15874: dout = 12'h000;
			15875: dout = 12'h000;
			15876: dout = 12'h000;
			15877: dout = 12'h000;
			15878: dout = 12'h000;
			15879: dout = 12'h000;
			15880: dout = 12'h000;
			15881: dout = 12'h000;
			15882: dout = 12'h000;
			15883: dout = 12'h000;
			15884: dout = 12'h000;
			15885: dout = 12'h000;
			15886: dout = 12'h000;
			15887: dout = 12'h000;
			15888: dout = 12'h000;
			15889: dout = 12'h000;
			15890: dout = 12'h000;
			15891: dout = 12'h000;
			15892: dout = 12'h000;
			15893: dout = 12'h000;
			15894: dout = 12'h000;
			15895: dout = 12'h000;
			15896: dout = 12'h000;
			15897: dout = 12'h000;
			15898: dout = 12'h000;
			15899: dout = 12'h000;
			15900: dout = 12'h000;
			15901: dout = 12'h000;
			15902: dout = 12'h000;
			15903: dout = 12'h000;
			15904: dout = 12'h000;
			15905: dout = 12'h000;
			15906: dout = 12'h000;
			15907: dout = 12'h000;
			15908: dout = 12'h000;
			15909: dout = 12'h000;
			15910: dout = 12'h000;
			15911: dout = 12'h000;
			15912: dout = 12'h000;
			15913: dout = 12'h000;
			15914: dout = 12'h000;
			15915: dout = 12'h000;
			15916: dout = 12'h000;
			15917: dout = 12'h000;
			15918: dout = 12'h111;
			15919: dout = 12'h000;
			15920: dout = 12'h000;
			15921: dout = 12'h000;
			15922: dout = 12'h000;
			15923: dout = 12'h000;
			15924: dout = 12'h111;
			15925: dout = 12'h000;
			15926: dout = 12'h000;
			15927: dout = 12'h000;
			15928: dout = 12'h000;
			15929: dout = 12'h000;
			15930: dout = 12'h000;
			15931: dout = 12'h000;
			15932: dout = 12'h000;
			15933: dout = 12'h000;
			15934: dout = 12'h000;
			15935: dout = 12'h000;
			15936: dout = 12'h000;
			15937: dout = 12'h000;
			15938: dout = 12'h000;
			15939: dout = 12'h000;
			15940: dout = 12'h000;
			15941: dout = 12'h000;
			15942: dout = 12'h000;
			15943: dout = 12'h000;
			15944: dout = 12'h000;
			15945: dout = 12'h000;
			15946: dout = 12'h000;
			15947: dout = 12'h000;
			15948: dout = 12'h000;
			15949: dout = 12'h000;
			15950: dout = 12'h000;
			15951: dout = 12'h000;
			15952: dout = 12'h000;
			15953: dout = 12'h000;
			15954: dout = 12'h000;
			15955: dout = 12'h000;
			15956: dout = 12'h000;
			15957: dout = 12'h000;
			15958: dout = 12'h000;
			15959: dout = 12'h000;
			15960: dout = 12'h000;
			15961: dout = 12'h000;
			15962: dout = 12'h000;
			15963: dout = 12'h000;
			15964: dout = 12'h000;
			15965: dout = 12'h000;
			15966: dout = 12'h000;
			15967: dout = 12'h000;
			15968: dout = 12'h000;
			15969: dout = 12'h000;

			default: dout = 0;
		endcase
	end
endmodule